`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EeIOalsB9A7gyFzgjBZExeIPJuRpFELHlfpU3L/uqPMoO6TuIez2KobOfgsxw4FitpHwSA97/lIN
csNqzUP09g==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hwzf6tFLlGdH/LlAouRRMzleWlGs8Tvfr64AeA2s2z4reQzhfo3uL+7NKshrdnE3tMEN66HYuwVd
9xQlnCboKstjE9oTcxVT1Q9+i6ynCWa3yDpjnUvWm0p5bbxLnANX37Tx0FTTAfpo8DSKKm9W9UkH
5GCk1+VjPB9HCpd9nRE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bL2EnncrNSLn2ffq1uLRkntupOO+jbrSmLJY+5LxOcioiLBdds86PhRnmpvnUOMHuvC456xH0laA
GUJu8mYWsLkeJ/gjFzllQcWIPJ8fmH+TDnW5/yyAde/a0JpR0BbhVMzIYr60Z0Rs9B0t212q0Gi5
cfOdS9LTaW5pBjCKt0jNfdZ8Lr4AQUDsXpboqkvDmK3/+QJqqF7qvFtia5MvW70KQywr5vkgRws1
BASbR4GzizLUz3PzW0ZpTpLs/v+rps64Cwqc+09rCJXCFOqMTOnvf26vB8oglq7BMh6zBeWRxEuP
co0bzIox5OWgSFlu3oTH0cogMWKub8qQURYsWA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cIw/9EXCGVcaeoMMOWuYgFWlA9RUYNad2DCpvqx230raBxPvQNhdOwE34j858OOUuWrDVHLj1nWJ
y5EJbcyT1Tah86TN1vYqo8sqn5YXS+1zRWIej0AYDEi19T5qjqQjxcf11goih0I+aTjhgw55UIbx
DOlEcwyPrQQ1bBWTza7LH/J9VH+m0Nj/ooSJpuXCu3H7BNulUXfTKVRWBHnUEaUIRnumtCzfbcC9
ERqZzs4FrgS6flY1m9XbUdMT4p1Eo893HLMAHq10sTH6EHY/8n0KLkE0TdZ534HUCGr6KkB4RIDF
99mj7IvY4KQjySVBm3SLkgpins9y6UuDnCijkQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IcyVbDfeKPQ4Wv8Ubt7+Je8EyB4He+T9m7hctmPOEOS01haLEIPmxZJ+0X54mZvQdvPqdj7E23u1
R3OAzZqlLWLW+d0PIGnEownI+S9ocJwuizHj1sJuwEI4jfxmJNZjE4H7mK9ZjmgjaH4o48SdhJi2
yTDL4y4yJ9WH40IPNyPODb7zhqRTxClMXzjuJVpcO9fl61K8ntq/eG0XNZEJOUgYAk+JXVhPJ/R8
LP1drMB6yJI5AgR28Irm3VsSjJoMYUTX0eURD1i60OoVxl2DyucunlM5CIRZ9EHKoz5SjCNfLkmU
FtKjFd9bGHkZXD09XWdopli+1qzB7QvkJwZtJA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ApmmzO+E6sydVLZl1/2U7QnosCNZyxTsKqLSJRPek46QkWcHHZkNFVIHCIci4gSId93OhQssVzwz
WXxP3kwkA1nXIZbFYCJMBa9u+RSxeQycrHAglmUYWkuVydXtuVb2yoM2k+rwZmSZ4EL9o6DJBzpF
8rAtNuDZO+/14GwY/z8=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mLieXakPF5k1udgyxKQoGQOFSmNMp9LBLBSpMy1hh3mZegEUQzRC/x5AREnUXKCJVi2A45mQS+/v
sWYfEz/mEcmJNfzQRumZAzzIhT6OZ1BKHYHb35ddARKqGfi1VsbWUgVRiujIoWzcq/UVTRYREjX4
QTMnCGRVa9CTZ5zSpFRgcb6v/R9mln69hqjdTg41euhxw8cfIA1i23jDHJi3nWhqoyUvQDcLM9/8
Dyyt1tIBHV0Mj2Wh0eMPypOfqhIduKFcpK/XdxKtvUexe1DxPTzpolzVZLafUNx2epnjraWTb5kB
0Z5dogCBc3Gek9KtkaoCoZYrz7kpzUy4L2reXA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 129920)
`protect data_block
Madrr6DhWrslCyKqFPC3z4siET93RT9yTmQA68P75h6CcF6lpZ15vnUkVtl2n4cTIDIyldT2Ue1+
7KwKx6sgjQzdbuoUaWfzlEqFqPeOQWaZNYQdS7WQ5u0Og93RQQ4LxLn2inl6qs4D204C3RxXBMby
g3bYfav3BwJlDd4b+6xPo3pRllD9zFFxIe5Uwr+p03pUhHGNI3BgDYgXAgMxh99dGrnmdtFlVFKg
ckcsiCeBncFBuQQnOQzwn7hAj3unf3xFoCYj9rbGUj1n7TT/lP7u/ixa7vNz+/dXFU7oo8zKHkHV
6/veVyhizYgfTw/BQQblUQwo3SexxKayS7wIhMH5VnkpaSiiPpmriBojkc1NmLUwuipgR5t2vI/i
lPGptjeDI8PWI6MMYUX+vN9AUs9wu+a7UDTLAzT+nBautQbu/6HKrZME+ldgwYqDcpigD8BIhX+W
tzL8vzxfAA6yGLzCO1tVuAb20Fm0xoDRCebSND+CzknNz/+zcwGx6RWaI6KJA3gsejpqCf8E6qEA
Uc2ZL5JNn032RTC6HlTeCBYn8wM1bHiNB9nyRR8KUp6rkal5Xe8eF2Nkzp9TS+LJFArxubrCTFDI
c9BcYeR+ArCMjXZoKC+wKRVSotGQUUAYT0XUxPCfFBSrpxsFICzxVVMpPG5M+15RMbmI3UL5lQLZ
oXUzSVLZWL84o9dTgHhYzuH7S7hLbthUwQsV7ibPBqxjissYamqN+rdAv6qb1Bq0KDqutaUi1ZeX
kFQYFhR1wTQRip8XOZXQLIVa+mOVTOlbpkmtj6IAj6YACXAdXQdOKuuvocEgDjVFgZdsHWR7oDsc
WCIv2AanhLRZo4CK4Hzzn5MHPW8xSx4IJt6cCprQmPAyb7VBjwNUGGAVi9qjAHoCSylFwE0Dq1B+
VLhiQHrbgwmlMJe8zsBDLRoHSxJI5oTX6R3rMnekmmtQgoy1fmogvIySSJ99gC0nwUPesSQ9jnRq
FamXDyvEtLTFWRk9YaXpsVKliHf7X/VW03DhWINIxe+XR/HA/eREV42S7yRAzVJr9icvPCoNR1K9
PgHx3+aXP6KngemTtZnn2HLW8NAB/3ZQcnkQ2TNYq9PPbziToEDTyNfWIt80+wvGze8R5bFsao2F
y4daATwYpMmU7hZtEisJWmoVHv9ZnZD0EskJwxqbw1KWvApmEUjLKCuQLX1H02yXh2McLXkj0sWH
35dqT5liJnwRIE6GQLfFtjQ+BVYPrF6pW9EfTy03+9tXdcx8S/0Yf77GYEkk38Qn0yfalYJ+61ej
2G+8FVmarlRC8f4iKnOvpNnSV2soeNi2BuRSrQJQrrnVnC4JjR4xl8TQ6j8cKfCBydIcGSgD7idN
O2YrgPwmRE/gYMig8OCvNKt+7CpdI+mnfYFfj6lGxB/gjcGcrUnwnRHtaujyv3W8JT/9ErpUV5QX
zuf11RuQ6aHKst1LhB1zLMwoxvIfg41FAwXcjzQfu0Gwm5L4fKUbA+DZld/l/k1yVuzRAJn32iSz
7XjJeNDB4eWrofvztp+mXOTblU/e9wo9S/ucVXHmG9NWIdMhcIf4ogO6ovwVcOcKaiMN4u4Yuwxy
mGPSn+6YH+CdKTfPpCk0ZjDRPma2fybnHW3Ui5Q1LnCz/B9YTetCVNE4OklNudTH0Y1GuI1owGbd
H/JwqBNXfGMDNzWBmx801KAZj4Kx/p8pD7ZXPYAZciRpZ1b6VdJ/2Vs+ts7XGsqBewEd4J6GbXMO
uMQFy9wZIRQbK4KZ3V0muLrt90uu7yb9uZe7vKK9x1olZUZOEz3jgC9k+QbnxpBs9w82VFQoEHTS
BX8zytzxBGqJes9lELP3CmHqB6EfkDD3+YpeXng44m5PluBd+K3lProSzNAUKAVBqhfCpuBFTSAx
wcFE6bB5VahJWy0bjbUnUPfHbCv35BnhDhzXReUCbiBl9vgxOKLOufWsPg1Opnyz4Zfz5RxRcoQO
ROfpwNM8tUNwX5FxnTBrY5KhSSy8mnApNkfxNFnsmaU2RRS/aWvaUvO4aiMKu3MW3JCYIv8ZfIqW
9VVBOz9KUfLlaaNtJhqC4+EwRSSM5rYijL65re69uIEcuF8rmuEvYTBw+pnW/w+uQx9pxmcl/J4r
6lg1o6w83cAGTkcgGetnrADJjwsgj20n7BK+f+8OcnbOy0Nvy/53Ke29S0Sl+HUoXw+l8/xxN9Ii
edzkM2ONLIBg09RoVJ5OfH/eEx75NltZRBa3UphY0fyoqmvSonct6W5wgTqLfItoyYLmq1x0X9fK
EA28fYPgAmz4jADZrcTFG6zEL69gJ1/hKSr5nPag7pfV+GrMcWwX26F8C2NfgrEpVi3DWSf9+/+n
N6nxZ4tqIr1+d68eZfKKN78XR2eBUYPCaUYqx1l5sCI3zk67YSzvhFop07ld51TMb67UN2pVelQg
xM8aqx5aam4R5lx7ZOLi85zZc2RJCeQBt1WEIeSVh7UoFigIc75bnvbbxWhGq2gWHcAkLha1Y2T7
VtfmHdtZKcrC0jENsOzk7DmqA5SRzx8r0/dMJcmmm3OcbNLiOIvQf65SyDyo9Lha2nOOIvTHXupx
uGog4XU/RXuQJDsYnm7fj/Rr8aYMVw6Y4dnNPooBkP7sZ019tKxm4T9lwsZBGKcSTOHnPYnn3jzf
j8qLDUqjg0ZgKeHR8U4wDspvMj2qurjNp4K1H2Z/G0p/gYUp6WalwKrNzhmOPawg/Hld8VTiYDEA
Mxfnzx2VLMNODcf2FdgxE6phgutnBa79u1iO0HUHFUqDqNPqt9D4/zURf8lywnk9rKTi6Rr04GE0
HTNPFGRBY4ANQpCbdyt8pzFenwbrqOC+2cctMUJbaCSgzl7VSy7LkL6rse+3wPrWg3HhKeyOxisc
GVfEKeu6+lsAv4lnkpgdArfrHgBPIz3ggxhWt9x9S6GDUEfNhMEhKg2ooFWLpW7kKteAbhgEy4tr
OmOZRKTlUUFwLbEHBKIohn4VEUjEAfaTD9b4KYACHuvKb9BgDNZklXx0KgGpK87YeAALJeqY7z56
0M/JJ1BalqixaCN3XMv769rAydvlPPK8S7czZ5eKJ+PLoz6HKvif/BeU72Xt2ZKfQzzt/WkrA4w+
VoB1SykKgXzJ7HH++o5B6HHkYPOlfmBQrvgnJQ1ANEN28L54yaIzrLUGXBcnbHIfaHIPT9qjo+lT
T3B0Snq44eRsOhqCXxbkj884Y+FWJDcUxAMWvouzrGR+BbDaDie2JfqdQ9IgRx8wdvkYyr1bzpKj
tiMym5L3ywFix6dMfTbzy7W1JljBXtf/cStFi3g02pF+pbOLsIEgwrvRuI8v4YKc1ITpnO4ZDY3f
IAzg49542Dy4nSCEwJVAGbTxvmBduL3UlUR6fBQi7JXHE6cozFdbj+SUgAwvXnD33RarqGlrYuwU
UcsucfMTNkltIBd1Mm4/k+S5Bc0jQ0417c+wasiIwXWv2zXD0GZ4hCVhgB7XHXylBErv8JkwKlrz
OBPAUN+J6E5KC5bqWIUQWnwrJrOLTSggITqcE51x161uh3Gwvjz/tvXq6njWy+Hbs6wp0HcDBVi4
4L8hJp2dXmt7hK4//XV8F/nyHd4Z1tuYu4wrnwQziQ2E1fVHcXuwPeOq4QfuarmHK/TLsDppmDGc
F0IHe1spq1o8cCLIwhVZ0oKdIOMQYx0N3dE0iAwQEsWyUaVhSIFnbkMwy1mxihjeAdY18iDyZq90
fM8MXHLekvhHZu75tz5JjlZbYgaMvoMtBwEhMGICONi1/M/HZmfFZJjx9wuF/wlE313cvqxTAcAt
LVVbYa7qBRo7tvcfrri1zslsvKqnZVF5/52Qegz5Sq9prXqcjMa8Agf+oqK9pAligxkqO4SPZqDD
UgO/VmimomncH2aFZ609eFjrUHosnh/3ex1cXHOI2U4tKAPr07yusREU6JJkL8JbeDXeQ4M95vUT
BG9VT3dJSwmxZiFCyU4+rcBr76ambWu1YGE4h0BunYbVbUHQJWqFl512+K4NJ2b+iWOj5Mu6EAu+
VZGHUae2pO0Xc02wosEw3v4HmCNY553YbDtH4pcrjONJESQyZEkFF8N0Ymre5NV28lvkqA6hJwnN
egYXr6zcm4yPlACeoPNvpere7TV1YRbjuf4oAkA7UpTeHcUrIK69YxmOhtfAMFD695m/I3WThoV1
NIMixBSl3gaI3vW/kn2H3vbNL24wy5Ge2QnkYcb4xOQkb2eyY7Kg7OLacIRhjYH+mR8UQWgHTu6/
kGUIYVES9oqKr/1YbhqFmEsas5aPmTl2iTqoryFGwM2bX8mRiYw2zPDUX/X92UI6Y/y4+cRVt8yV
bt6dYkfczfql6v34krWQ5GSmRJqi57KImvwE+TWq/N6w32jad1XC+b2RqGcQVgU+DtS8WNOgmxgz
2vg8m9v5d4T1pKXhB2bNwsXQ49jkYZEEoBL28PIz4tAKMnbcsWiymRSZSyqTuq9qHojuGahCdp8L
CQCsr3oMCLNzd179V/xXG7dwkIN6y0y7M8hDdicEPgl+Scaeb3rdp2Ko/B5BOCXEy4gH14VQhoui
AYpwcwrC/NrWi16w07HZ1239Cs4q3mWhldMC0DWnGKj/RzALZLpEL+pEt1Q1+pMMpK1ATZvIqN7v
SPzweojZSIMywFYNklhZfEjVIQyxXbDVjL+uvfIU87HR9aptw2KAgmUTZWuAHpM7ePft4NegE+ZV
enkIdsjBLGN+UeP3XoQW2uTUi/kk0MOKa4Lt+ZiFN0sJlQRdOQfFf21O4sEi0+szIUWlehGg+Dag
mrvTgqkN8DJhNF9WoyiBU7x8qvdI1m3l2+PfnDyIlJtTv63WlrP+0EbJ6R/2MVZU/1nmW5WCwPap
HSQ4RWQqOdjWvxAMxK3endb2i0jBhRBI4Le3CkTgbY/6KWXjIWvEIEGBchPLO1wro6mW/szVPa9w
mUd2SWMY8ald/c1NSxkFmb93NhDpBXMM+yCePFKZa0WHDmQfeMDz71AKwkWWHJ/PZbZBTZLc6H2e
U4jgR+AnjaHyFk6dmXQVBgTFCZs6O/GzCpcSIVdnIvlsAE2TO9i5EjI2r8fxriRaeK5D9JfoCGga
VOwUyqGpqHHwksC3ibr8gKIQU9a2w8tJ4zH6Qnm8AB7s67ZaZekG6SxiT2PviY+adLJZap/Rdxhn
Tae/VPYi6rp9ZF5BOmRy+Wefbfz0qdlO43QMW7Eto5X+8OP8CBKRB0XuiP1omf03j/JDVZ5Lbwbr
DbbgFbcqFXAHP2uupEPav6lGBJ7wbaImy6LC/UBWfX/wUG6biI36Fviu3u3B09HGj7mL5Q/p41E0
DXSxoldBVEurnNbry9uYz8Uo4vtU7175QOj7UunA0i+VS25c3B7l48RmACRZc/pzdU4bRMB2WYrq
JYPysNO4PwWMw2guophc9f38Nq+zITi9H4VzzDwCGOftMECQQyP3x3lItKWDuzoReVidwaBU9lbJ
CL/x79jA7758IFzjIoGI4POBJK63LFe8zNNYeZ9wspNm2giXAwhyJxAAxMZf7hMzzYEseOAKlOgx
5/6fUdEwfdVeRWMU/NFG6oLX8hjbwXnPNtMrbVXvAOl9QhNd4mGYHYa6uscXaviOZS+w/Oa8wFfk
Jp8ZlKrgZ/P5Trr2NtbP7ysCssye96rVuDM9YdvU5Xf+x00ksLrAxLSPPPoCFvdTHiBNrJ4RnaUh
RKf2BQAJnfaQRRzRB2F18QdaV9QxnMhFO9eDpyDxDx6RrvRIHrC+w98LkGLajeGXgJ/fAJRYFl24
Cajh6ne3eW0xBeeG0QcCYZByTGL0iD7egVecilvGYVSfqys5la08nS4rPchj8k8yPKiyMsi+zmPa
OWc1ufrUyf8lxeGi72ROIx0h4VdMk/qPtbv8pNMyNi8q3lZfNsaNNqakZfD0PYR0+kJh1nDPGxSF
4UVipquoZmfla3iuInYrStz/mbmRik4rtrqggaS1GcOJaVjDIJqESHWmPlyCHi7O36mE90CwCPR5
G8zJpMvTAc1E1IuL23fXdSU0FOE0vdEi0FkZPX5TSfc9gAq6Dw20epK7vEtXnqIjuvCBizOnBHst
80uELJA/K05lFEA1gyKshuqJNlFZ5Jwn78Sbl6lSTJ641f6KA/EnbIVDtvCc7Y+3tCorrSSEWcH1
cPDtPbBGCsU/sTbfFAb+xgATGkUiw6+4HAlsatzIWbBO2ZWVmBBlbKRT3aJ2velHJx4TLxpUbz91
18h+d4YlfrL6c+kljXsAwwRDd3ec716NBHUeu1pjOSynjCDeTl+sZ1j7wX9D8ITZ6oz4Z0UjpXHC
2+Wa2WRIoYPeYd4fLVq7hFVe3o/UiZbmcvr21s532rOZl4gZBrtbESnXCahpi0n0Y7qAdbmou/cO
zV3XlKh4LxC68Fd100jDW264poEmbrs3Y7hRzF8xS2gMIL6pyreJuOxcv0uJ3SVDLng+mB73dSQ3
KSODEXK2U/duCZQ5MNz3yK54AkHKtJ+KWQUKKZB+zmd/TsbLX3fqblDhjUhibmx6iYEuoXt+yYtO
2hY5nq/UnlN3kVMv+SVvuGdpF89e3/rWeOUXTBcF11T6dGDeFwtYqL9f8QTPRdqWi/YPo8TCm8pb
JTayYMEFsyn1TmaQ+cPnl94EcfZ+OFn6bEPAIIMmCuYGr6QSUEOUVWGawCfHrJVyahDF63rEqQ/j
SIk7ouzdf/D6c2hEa1FbVtgsBo9NIOdRfYBd9/kp9aN0Kz4rYYn6Pc5+TiwOlNSAv/NVgwUmV1iL
44ZC3oglzx1IRDKE41nTG0o1MXM0xomgajK8yk4XXH/Wi4tf/IcrgLNCmmRC3iDEpb7AJ1U5IB1y
VRr5NDFsHHSbmtZrzN7QmsOhuCb4BA1DT4bqyLe506So04Whs+qKP1jWx+NgUBH3EHiFSMzqncYk
iUXaElGV+WkvzZ7UhgtMfdAspmecANVPfaxrII6nTYrObfkh9L7fGScAo/FRM/xot8nCpNl12xk6
LfoM98Cm8CoSLW4roUNvJTc2UmZ8wT+4o1aiZANP0d9l0wNIpoH0TtosRnSj6CtbRQkRRHoZzJzc
fV2vGtTYLovcYwf2mkV3fVS3qIIhgEO5Dfq23MQOAdGeGCYqf6QbEiO1JDq+DCrWTrw0Yc4PallU
awiI0r47xwrtpy/wExe+yoz3AMUbhXosYOmMOGvOfA1hbnCjUOKgRogYeU0zQDN+Gc58oqaIt9MM
3VMv4ohYPMUVNjlzhcHDGsryqjUSa5oC/EihclDx2j52S2ViktL/+xO3CF5rkP6lN/qYXV+dz/Rk
GJz8nhUCcoK20XVgr5edyaA6GdGjMyKz3HU+HMLmNZ+65cGpwklh3ysGPfI3x3wa/eodObz6pFaC
ihXfvj5XOupVHJLui4eMADt1ryUH/EDmDndeD4zKxHTzTgDACLPftivPGOOZwSPYkPVSt6uoMoNo
NIJWZp67vqA9Ns5UjFNvrhJ2hCCyRa+RVYKHTWleAso9OaYtHsf9dpVrHfpWEDNX3mJE6BEGrmRS
AtS3P9ibXFmyPSHF8pGb5JHoqWZb/NCsU/o2SJ0GFeI8JIH6nmREKaBKYXx6LlrVtEwC3JEpGGoI
VVzOg40E6y6cnus3ofnbo01uP0PzCoMh3BxGfbii7hel2F2JjLmiz+Y0y5ym77M5+0Qw1VS3RRUb
pc4YM0wfDCDtiYTfOP8UQFg5txDKXtWAlg5KRy/u36Izl+QVztUHuavzhC+jAYu9807FbJSrssMm
QV3SUSGzUDHsyumQC8vH90YZixU4mTevMnDl+apBnATPQtRKDut+Am+y8coteRrABtpOlvW86jVY
iUDq9oAKV1hYiS2YACjVSFKRfPV3X58+MY3WcOvkNJIr0zqzWfM5yPRLDguR2FylluYmHv68rYe8
zCKJg/wlQMEI/eF+UYX/EMNAxWfocAiaLkbwbjpk9AKHOLu9bi4wYSAScjyK0Tykya2UbS6bD9mC
reL2w2pFR7bstn79K0w3nMnK/8HQwNxjqxqkRbUK7v0N4jIsO6q3mwUP2vz3PDPjPJEKGm/c4klf
OAgTVOKcACV6AzFnmgcGqzFcVC9wYsrIxaQ+uzroE2EQ7noNYRbj4uie18hi7o9v/jVqOzh0MaAY
16ouv5UQeZ4FJpVxfS/yZcrW5c95yoNDFJzSEONQ428ljgp/SYEWf2XiB82sxSzogMCrHtgVAsk2
ksV3c0zI/HunRXb5wcfzaKzpcaW9unDa27NmYoym+yPBVqV2maJQNMH2cqNZkLjGEjqC4lT2vMAQ
ejpJbPneIuOqYDAueXnf6PDbyZ8fdm1wFf1+GJ8QG8eEYhIl21iAktcOVQHHOlusfo43pgc86/i/
dsT2Lw4VBnaxQolK8/JX5otubvDbejak9021Rg/UjTsUHI5Xlbaj9/0TcM4mkQFVJ+HG4okk0/Zd
LmlA3UNLAvCpblkjsFBMIoPZ8iaYs76OMfNeFmudHJmoEkPOMNn47ES7KQTY8n0/yzAQNLn7Il5q
uuPSx5ZGsBObeVeWJ5QCnKXsYTkxF4prF6y56jsqw5hYBRLZllsr5N4QUIKV0DExIGoi/YgLm5d2
QEBZc62ipNvq+YgeeapYitZq8tXnP4kwVKFYIXft0M1wWjHtLH0xmSUV9uCLG9m9fiRWty2hstG+
/ux0WKANgSQBum7ohMmy0H5dUvnuyqbDHfwssW2n18yDC3x+GVRfa9CVVjf8vfXUuiSmVHOho8V8
Y++QTpktI3PA7Usy9Zhu218PZUEGgkg8aetNrZPO/dqyGlqE2NQddGYiKHCILcNkb+DKCu3fYT/3
5aEb/2IVLD3PDB7bLHgTsscHTttu60NmuMsq9uvbFLTmyzQYDrvBiD73/XDzW2ZwWKGCEpuVQ67I
oS3v7Y4grj4oIUZC14KsEhZPtmKX1MdnxJ/gW0YEz2niGKc2oNv3YD1nUsxFcDou6ZGUjFwY4mbm
FhsqFhbdAb+Ax3up4eYEL68ZWjx0DGdolW6YuXAQBZc/efk8wVOTlc7xqGEsKwTeQ/Dnz4AjUzd0
QSQ8O+9ny9iI/ViZ4lr6sz//4CcwiW+LuzHPcG0Cz4Azzh4TNXN9A2qbuI+DiiJI6vVXojNnqsTK
w+4bWfiicdwdhl850nNqpqcPY5pY3syBUWiGSr2ODXjjh8jmKyxnx/LdccS2XUwj2jkVc9fGyd3l
kQ8BwJ0jMcho5+uWb/8rmJWV+2gQSL6+jsS3l1fiFOIXUmMRkyal6mbT5cvIDbB8H+R/ksBjkaGA
eIVKj7q0skv5gRDMTpMiluY2qIR/6jTBtJ0Sv4LPFG4Z5cDPzQ/PwvtdtvBAi9LJQTQf+q3gFZug
fTOCUYeFSj0SEy3DdUXEzJKddWwUhIplW6v9Vol+A8oy1z9VwqMHEj8PJKeHV2iJml82xHAa/Mrc
q6M2kk4RLasKjqGHmdUkw4pxD2Qh/3g000Wq2HemvFx44smWDCups/jo3WKpARJnxTfjLU91Oiha
3M5BohOPf5F112mLf0vjr+/fo0bXQE3mbBk0GhM8EG3ZvHQfsSnrNEMeVjICLAd97WjKiVo2ItWR
lpfbnYN2Mon4Rv1q4JIgV92rFIQh6ULDzLJKKeRRGu0y+p+FLHdLeivzMCXFecWo8ByIkdV9PHIf
6RnMg2PueZfsMbv/5BH7RmYH2XR+a6X2q5tF9hDK6Cyyxe+Ky1juvodwsvGp2HihymTr1QuHYNgp
XuF0VSdTJteTKDJTPyB6leJ7v9jYi0/rjTgcw1/k7zLEjp5Dk7Q7Px4o7P4WUg6cYPpjWfMP9ssv
66hIMj3t19ntnwOG9KTKqwz5Jo9UB4Kx9+yOQOd/fPBj4rSnCbFbGZdZ0FGh9ZxCnbATh0mDYB0g
8g/0/cVBhpgVsUEfgp5a1np6hiHflq2AZp2zSpsK74sGp/f3nD/+KJA4UYT2ZOrR8Io4FlXE/nUG
mnARpNCAMvxaDm+nyHUll1OZX99/z0Cj/xVbpBCv8MUyADzAdomfP7ClMz+HskitfuRxV4GVQwfH
tbG3HJSFw+VoZe5hYYEcn7ml5BbbyTlYFgt4ddya2dEKvLhtFju9xRooTAcwZN0fuHK6bqhoB001
Z+8KBgmpTcR3NTw+LKQRJsrEQpd8B5kRFoox3ONlvV7xy00PdppXGoIGd5/3CEuunosTPgKCk1R4
tNVinbUQV8jhylNOjq1/E6W3tWnp71e8sVQYMtks+ptlN4vm040u8tkvMmjMNKNBHOpT8FjRTyXl
ZPGCQ/Rbo3P+8GNpiTxv4oGfmASEtxuzHZwe88x91MmErvcUDz6pIAM6ikfAiFrx1xAHpJGY7aeX
BJwpKXPIj0u0lwR2sWmELK+agstrL+GcEPK3s0DhwJlzaPHDFYTzt0mQLW/c51qRMmsh/aNz4Wli
V4E6BpSXEGQEk367bAD7vXSqEMlamL2Q1YRLdSkNPE0vHnyYqyQGDiP8lCryM2EGEZsoDYVjKOTB
jv9iB3P5u7all6Y2SbbfXE/sX+TrGIz4/O4WPWMvEaO2hI4LqetcVhD0QjyGuVOWBMTjbE4R9URe
czqB//vZeMjOR/74xVQJld4OMLYyrV+LqMjCYAikqgpnEs76rAnLcTKrzTcyoqLJWSPy6yptm/W1
tb/ENq4kV+A/t44nMkeO1Ry01N7wBF2VkNvv9dhqQBR0ufcorJEOVALDu7a1XFkV58RgvELCwk2B
GgIARFbe/5WsKMl2r/hLy30sItm7QVStM+V1XfBJuE6YCdB+47KMjTU6vEB0OqMLMngNb4XLZsA4
3n7orGqiNFO52Woe56VSMHDV1GzWfV8dBHvEH7e4yvikDb5dFQ7aoqsUZprhZfYP6PcIEnGikk3l
g9OAEqB8xTq4/ruF64cTX37qZ8D7P+n7Cx5O6OrHny1zbH2OdEH6zYIPFa/AmHByxibULhBjAIJz
wbLz6UZmhbIhzGd18gmhy1hS4ZLB+FLUcJ2uT7j8MB2FsM30MXISbdBCTov7NlToOv/88E+t3A07
QJTSYT+EoXOLEvAFqD79OVHe10QVDRwzYxk4lsjJcOmOjQY8iIcJgAQHqZzvVTT3XdkBoF+k5BI0
jhzdm5qptH2BUi8X2A2CZKT4bQ1PDaTaz3wvK01nLWs/hCsR5yJJV5IDEqwJACOK+ptsfGVTN69G
xmwzVqqWdfhv+ZVqgxJqKqK7t0qhpvjvwTqVN70et0NzH0oy/2wsKaM+Aq9SkTneet6k/u31aGU0
40mOIoBCUS0oBzOqWyd+MYNw223ui4Rn+ni6G/4GZz1uY11NTOrl4K3U6TC+V/pNtPuvOijL4pIi
6RRuFbI7jTLXefpSmiRv8zlxFpaKAiY164QY+I9f8OYsuU4fAVdmAr+eijt6kuyH90dA3uMNmczS
OznihSsoAqp27CQEqtz+QPWufPH63JcNEtuSBe+BOdVqagrSJbgpMuUu7WfLnApxgClH+Zx3Ilc9
1WlSDJMAACOdBMb/+XdvtiTJY644Qy/Atu+jKpt6YocJxYDjIZTTbN7d4LOBl0kHyBiBcbOIFADb
AiUDByFvSj/KysxW5ruKsXBziqlkscLZsFtpzeCCR8OhyyMfFzTcJxAmVj+Wg97MC5HivnBntHVz
Umos3Q9H8bEy1fqI3KeL7uDJdxSXYWU/sM99gU1AA9gpDXxQCgmQFrtdesmF55DuafOyUS9qvC9e
YNsZcTZkf3UibzHU0iNhpF5PmXO+lE5XjVUBByiQ1BC+EaqAaHiHPrVOUC8eHI/C4uTMfi2PNhxX
A6bz2m2X6QmQMvRAhH2oDVK57iw7yesVvnDMsC4/SjsVklQeZKA4AakatWZF+PhNzmFLroipqHv3
LfKdK/bVvO+oGYPNkLyLoG8Xeq3YAz8vNs4RTX7Xng6M9tz5lWvnqa+fG3w1IkwIiQNDQ7B3Jvv/
Re10+9C2AAj7WXO0E/FD3W/YA45ItktmhdieDW4GlzjRipaph7XrIb4F7StF4VPrViBR43YAdvvg
oi04MkZJ2h0u/CppXULY7K7NhECJ2w/VzZmTNuSCTLlM3zW6tNKNXhcFhmZz9qtyhz7SH6jvkDWb
aXvFgHByg18uXlQpfPzvhr14Cyz4cG6nyBx8gs7DWkm8VWdKt6haUHNOdZw01lXlRGKQlQbA+iP6
UTUG4P2b1YL1bD8CduvLN7ojbMLjBu8yrPQXZDHNYGl2A8oDq9sXzVhABp5TgoDIHxsxY3EwUu35
8IjIysFSxviFEsV7VfMkDxKIacG0Kul6UavCo+3Ktl6AL2bU6zCbCI6zyTSq3ZSIN1l0rBpB7m19
hvzrLshS8do/IntL1WqaHrZtLOaNsfHyREp4sj3fJF+CCVCMaOvW6JDR4sfIFaE1nmbrJtyBoRJK
+oASi8UETFGc1O/xxfAXteOIH5z/S15KCKHPpofjjD69KaHvZ0bJB2+xGJzgl3cRrWoHBiiJvbu8
s0iqcmDlX4iXChkrQWUIvDTeSrwim3PXhoNDjR1KEwAWmp8Kn9xIEg/Thtm4wSOET0J8LoBZJHys
94NVWGdOO/oOtC7X8c9ZCGrBh4Flyl30iirWJ6+mJP06FV5F+s0qMMsgm+NOQVnPZTKKU8Kj55vC
SMhLBMLxtC8K92YSnz36A6iv1AWaj/tP8OpHGB5zPyIfofnqcoa9DMkvTmOTmKqha4WQYaKksTG0
iLLNzjsba6muEBQrQN2OISJPxAHGNKOJQ4PEmJ5awrF1Tn66wUwfgaq4neyDc4OXretr3ZXK9BVM
sIIgNRiIShevh7QuBFyFO91s6/KFHwpZ1k+hjx+MaoiNtFjiW4oMV8dEblHIbmJVqtpkI/UlZEpX
1Q7YMqcsp0CmIlKcW17EQwdw/gAMZ5asm2CNk8wFqwH/4z4dFR350dih+dNJS5aBnRiYMhcuqDAz
F9bF4w2ZsuKHaWUh2CJyD4l/VsA34MSEctd+xj1VV2gCZUHlsZ7BLmKsDAFrinCo1p30v8IoXqoC
ezSE4tSnn2r44LA7yqU4esh6WIZZQ/wdpyEN4Y+N+B4FPDI9TTTVYkVsgy8MaZMq7fyQ20Vcbhtp
zeok8Ti5cxrqrfVmcj/xzikV7MSwcLZZ4CuupM8vw8KsCqZ9NDCQwfUaDSaDwigLtaZIDs3OjEx3
nzyvmdgS6aTeBEXPSVTtqOy09xYnNOqxqxcDZBUHTaGjeRc2hZLysUYDFyML5cw3x0sdbc77k0No
EOkPfeQblXbbgZfYDN5DNdP059EGjWZIPdyi2WxFCUicbE2MKaUyVQgbgKx4052KJg05kYoAcLA/
cfLZ7oMWNmX3hZIYxXhQkrRLVXJZ+T1o5uUtSrHeAzZgP/S1r3qMjyBhQVT/5vZ9yUBQTg3Lgkbk
PD81LiJFEy366yc+dA7Fr0U8Rx3nWNz4/OYSWN/sH5tzH0G//Ke26Dl540CgaMM5o97qmZJWsJ2y
50iQpxuWT4BGMU3lZXSSbI4NpZZNrFzQVZWT91NvLIMdX74d16lzAmMb2lPFz8mEaIoR1Msrsqv4
ifjtz5luvpPIrnczqTA7ricQvLRRboxJq07nQVAo9TnjjeuIrbAbsf1fjlJY/WHaZ94t12/he6Kg
le2O947ASn2KbYCrepcdNgvSIUucT5DBpCR0aawVOQLFoB0z+3y2gvjnIKLJcngqPYBu8ygUReqW
WKFZsm/0p4osP/UhScCuNr/Yufw7YjfV3W7ZnpmeYGpeYm37eu8wufUsmX0vOLJIzc1ayNDB8zIU
z9QoYqtvPCTcsEvjwKDYJyz4wrkaifEYj5jebNCEwC0I7egfgnaWo8S6dzDb8pS2roAwGSJu964I
DoMh54AtcvwoSGIq/rfy8HlsEcIHY4kODpAoVmpkgACvMfmS1xq78hB4xgX5HWpQ3R95AoLqUN0i
dINGWCMb3nEJGipsCfAJmUU0dwIreBh7QeaXEECbF26Aa/xsGGJvsthQwsvc8BhrWLAqoOK0gOco
NkScQAadV60ygFXQbUB5h2wen4CJDFfOPn50XuswqypJ3ywLFLwbXzxRWuw7Y2WFfcgSsoxPc6aH
TzANpOtsULydht1Wa3sDICc72Rg38h/2VLZDCb8b5FJnB9zdhEf4RLcYR1nopoAkveRH7R/6dmts
FqeIc/zGu6FuwB4u+zfpdVhPWuOXYWoC6phSNIZjSYISALW/46A3dGaagU1xtxaskxikvMQGvWPG
qkRyrR5tCT8Sg0oV34JzlLkKpDKSGTcSjBDI5DcIMPFrGcfDAF+1+SH9qnAU/ttylDB7twc6pWsR
0KyeX33lA6GHlokWyCy5dr7KpwESwR4mdMPfzycJGLESQwdZbTxmAqQY4fp1VtClKddF2CfJCehk
ibyR78xLfRqn5omJZjt4udnBvIHC3F+REB37/bvDrrJJvXC9vM1aLhSf6kclTxJNqJvWq5Gb8oV5
00/EkuZITJN8SCrW8YFEl1iwv9CtKPm7hWd0M/4Dzf1AGG71VYIB2fflWxK0D8z2LKXmhyBVWb/Z
l67AD1DGuDolx1Y9rXtH9PyKYPpwjOeihTjybIeSIXDjcjQ+emAeI0yswkeoRcTrGeWbhSmLwlQQ
HV0hiDXL61gn+hMGkyllaEm9/u/VOJjYkZn8tLoM12b+mpSlfERiWLTHQjorGFlWfCYPC1Qkver3
L9+jN9nyFGrZkiQLhUi9HJuzvcGs4FUthWySVuWoRH6QLSTxzONQxcvMgv8ZyyW9Atjkuk06cJM7
Z3xnfBrII/EDVOcnCmYaVDH31amWhqDy8Eku4fGo49JGmTNzNMJwxEJzBbKHDtACxIU8udqUSh2X
Lhuocha91kwuXwB2iOx0CmLEhyZmJHzNKeL7tlJv+OvhIR4+fSlKJT9GDyQ9nAJ4SjLY+WWnzr8m
XVzN6/abjkf7c+buAHaO1ALAL5gMGyD2G+GofFkdpGf3GXf9tSDI43h0Z0Uwn/o+H3NdjHLfoTEg
ZB0qIIh3Jt3sNICq/b5dxPp3pLbpNMbgs0Z0xnR6ra0DXsUH4OvGj0iaLwffpAHYEJeTCAwqx47Y
QM0goRmAXuK/BU7OynR+Iky5apqUGWULlvK1f3F//kbDH+WIlIHjYE27pfO4Mg9Y3XCAfHpTQbkR
x2bRbjvFS5mhS9VEVwxPZNiwFTUN3AYQSM4qjY7PpCnvuKB2D+CDmApBQqcLAqyBrXInJOzVpFND
iXPvrRWQA37PsCpzyAwipIpRx6pFQmTZ8F9ySsPQcYlzgyhOOHPdax80JJuOihFxAyfHMztyPJYC
qHL2jNO0PzHaXkH7AqZqElhY1QxbXGmiso82tk9Z7ClB8lnhVGAFFnCKNKsaguReF3noKw3wymzS
xV3to/dxvvyvUPu/AZDIACCfcaWZ64zTv7F+3xo5nT18D9Gj6dnb+iE1g8nb7CwWNPlIMGE9GaxX
DoDuBhTxCjc8C1sSR174Wue/RzkL004TXo72EWuVfGY1SPEDAbhaaEemCzf/+Lf0eQBg38LGAdpU
0Dh8jSEXAh8pTQpKsRrmrmbKR9YKv+aZKtdx7gTO/uNWAWcZkRlMiNyq52QyyH8HotzLxBl0ZL3L
TnIVdRqlw9hHr49zqnDIyrXvwOmBASWj2vad5GW4PWps0Ka1gdA6BNvRlXC3QCVp1/zEmVpdVBQE
AlBrX3XFSb0scaPejPnfgTpJUi2/ChgNNyfCT1FtJQ2lldhp/Zf3TPs8SPh1aHNkgqnPleyMPalZ
Xex/0ngjXIEMi/7HZI28J4lOf6GdmI+RCHEbEqJYSZ7NEUN4Xo0vnrMqPTUasVABlZrNe0ja80b/
KyNWS7YsjFhnmrISFyHM3Ag4m8bMfk7zfT8SGw0adZCY0vJ1RtUaYmZmlXPhYAGF0cud9cBh3LaR
NWZJTs1/Cy0rheRMb130M9o/hTS1fezkwX2pxDtHPEsQ8/cRZWKcwyJP5U0uupLp8fNcclezpjWn
1seTaUFTdj1vFOOERd77yYzjbjIJQkI5sHKNq5v4IqtRMr1p6cWNtIgwg6S36zDhn8lZ7y5iAEaR
EdQD31REz+y+fRY1L5/RscLhYHnumdHgG8QFDWwY0yJ8WCWoZktNDi59V+zF4dfLxYHGcwnRwEAo
sdzuTi90qLO+fvrd0dg5GjykjZSTj51QycLzpeZUWp1/Yu2cyHF2f1G9/XkWhj+mpYCSF60QFMl4
1MoOJCsUbA0WBu3V/l9hCHGzNnXRCeGm3N2OZMAiAuGtfLaKcswsS8+AZMxkKGGl26tMyGPULoab
3NgqbB8TwTJbKZLJL4mHb4DuqT51wTCmfZiGtwZ6B6tKpx/FsITPWWrKB4u/MdwMNgBUxcT6QEc4
Wvsg23AYcic8KRyc8Y9urXe2wHojWY59Hb9XkI2xMMa6dXrsLrd2p0aYSS3pVbzYman89fVlImEu
69JLbp/81vGyzTaxxcOZIVD1N6DqW52wYmIhslockRw30wNlvkS5hMYMRivXQpqTQLpwCn8x1/qm
zRY8HY+fcAjiHwIzoEVYAOiHkF4UXcQXXljNbXtFKiXjtKjxATl6EhcKp9oyU/DePNSFw21HlkH6
hYVQgE1lNB3yWGfdfnuTP4UFRS4sCXyHtuEcXrmPiYIa/7mRHxNcnfFTDcryHTCqPbtR7I9uKbpe
BHCuq86+bTo0mMIRkEkjZYzaJhCmGrF7xbrrcJ7uUMyR1qqE73aTUkn0m6gHO/GFeJSL0jcsBGxT
icgfd4Uu9+9LrxAM0Ie4hKMxZ5nKS15sSoZ6RNncph3cRa6BG/8C8q/ylomkpcxJJlnZWYryGM3D
O4+CzIWTjHlHZaRE0kb1W8q5swflWgpE8aJMAEd+ZABDoi05yVr3Lc7iDzA4o+KWUBtKLA5yNizQ
cJrX5v7o+D5GERZuh1pyKalaOHOudlQaBy39U+7NpR0b4/d1kQb0gl302axv3TZHJ5LcYq6Y1r6i
5urAa+5JUTcOF0fghlEW/gMKb+xM2tb/lUzNwwR6ZAfxFGDFgvt2txmkX/l0hcV8C4h5jBxI2tzL
5IVb/JiabwJ+/pRyHkMquLdVi705a4z1F60jGPBlA6fEggXI5K25EcJc9AzjDf0zWEogsbS05C02
8jL9RxulVIhoGvkmgUPsitePAzuo9WK+UB10SxsGjcewWQk34AsvdHNiB+4eoElhXCn+cuKredNY
qa0oiZeAGWEpN3iqboN/mEG5C7xi2qBEGy5qUFFQwZNVCiC0xPX9PNrtrFm00E917jBbRzkDNFWu
ExDFP5426PSwkaL4MQfox3Uz5BwdXcvn92RTIX6ylV3N3Ggr95EEpNhFT5ZWMumPLGed++alsZUP
872UTPV0bgS3iXkHXMslaJuf3lKGfvw1LVVYxIhXu4BsjuJ+fGupnC4Ksml9l0H+C1xdBWwjWKc/
cs6HRZdWxif3/6YfaCHaKYOXEq4jj6zPXGD3E6hr5RQVAt7PkaA7UB412i1wgNrVs4g/A3ejDFog
bYox1J+/f8Dhh02Z5/0FqZlqZcxiDneEOI171UF5DjJqOgFsY+RqH9qMATLvsD/m1Z8IA4Dg+AhG
xg1dsHVESbZDyjLOUr9Xg27WwabKwhIl32CIPCZCg2NfXXT8LdRf0bJNdzDUSw7ULATAzs9jVIrJ
J9HPWalq2GYuGZhSJtK789apYXxT88XQrRHyj2Zvyent3k84w36Jh/oivWMjt/22vSRN39Kr6xIv
EM90fAetYxS5Gy8SKN6ptwPz87YHA6faXgzTGp2gf4H6md26WDhF3B5gh9ttjWY2dSMnPHmNwbvo
AP8s69ncFvIhIkNXbM2jxEvf2KYPI1plzk5BXpsBd4Av8zREdmki6umbh1S+O83UijYqguwPxcHQ
/YwtLobSnufl7iTpthNYsRblYmarAfDV51gPU0o9/TnSPU+b4gx6BlSa4oVj1zFhlr6vwv3JnkH/
CNHcLB9+sGKVes+RJcRXkUYRpEAp+tqGCOFk5rUkBMogV1SjHN4GeXOEwH8In2rX1u+J2dPlAps3
diNwCuSJhEOfSrDiaJ9DhVIzy2nkZp+EGDE+5alH57mTW4++RF7fF2XiLOUR6eScXYrnVLcsd3Gt
wXORN54D6AqfWEMFy9z6GMAfM8vNE+QsT8m0a27aG5Yb20dF6pncr9xnX+4/jyiUBabzcMVV4ZuH
GXx8REv/SNqZ4nBtLVEv+rKKUU0PngBz7JrVC4BVfzh9x0K8DSGPZU83yR6MDCqKtv5ee5P5qAT7
JsF1CNHOiABObcWHGXQKeRO71PvIN13iSnXMRpFZijEOo0d1cZoDhxVtNfVG77VzFKNLQAnn2zN0
ngVm/05zB3Sgh3nL4BhjvnoMGtIOh9YUR8mrgxrx8Wg9dFd2f6antNtmXWByVz7SioEea5MVLub1
HhRqW5neHuoGrV+hv7J2PAGJPSdwedLhSjhzuuI7s8iOS8ovKaR6VTiXxn9sK6QHhE4oa91H0DPs
P+DwZKlnWtgGhUXf7olHfS6oknRKDfwL6pK1gTWGgd7R8k5krIANBunde84GpolzyAA+1J7qAZFx
LufgApEsO2XMYGumMp5wOVw6hiR9HhIfb3wR944It795RYSRuQ+Xu690aIyIydMVC84X3rE4sF0V
N5HPadgy8027GB83DqKSziZzaqkkCzdoFeDeznhTZ3XexjqplrOZBZ8kO21XnLrCGwYmZ/9kklLA
iCHMS7tB0dHtK+kNsnAZWxqVm6FxeqLTV7r0vT4cnJYjnj2jilaRSQ1TdrGaE0M7y+8twQU1Unu7
teTNkJ+d9EYqgnBoZfyOWKZ3etEBqWr5oZFfnemX0T5w6F07Ccnf42OoWvgHzZ1GJC2zf72Vr30N
kepH5JIP77MZvma1W3+D9opHLA3iWqH/iQD4phwJY+vDQbuTJ7iY/RgtEwxz9clcqKdFCPW8AhvS
XFRnKTli+oT/wr608WCXh9obuVNvX5ssbqX8AVobw4woU+QgA0DtVZZi6LD6dGoezmF5aVT6hJbV
uC/ezpRDVJ+Q4g3l/q7GGH87qM9oGpABcRDmHTjaCC5AspZv+FhbZSJPS8kqMXl0g0uuuOAan7uX
WDyv0B3MSExFcD85YKkfrABOKuKb14SgkC+mxc8hviziPKaqTxAn3rBqK7S3cbHcuMMqRCzTtjiB
D9BwNQn807xwz8JnzFfqedFKezEkToaerSYFRRT38phEzmtFAr2KViRlUNlnk1AE22zSpjjLIRmR
MOPq9Y9Uvqr1c06l0NxvnPJvSG+bE432lxoHCKP1K4mEiXnhGX6H6yWiS73j94awhZMf7WGvumYz
n5Lg/KyWDJ7u+Gp1h0+cgnYQHMW5hfn/1JzU0M9iEaDeAWW8VJMcm3DPSkm8xQZxlmL6KtNYwAMs
M0JaZHWXGv1tgWsQAwInJCR6E+OZuhlKEPGd0a33/bn7q//+PRozZzLdNHp13LfeC7H+1+3tS4FQ
C2H/cPHThOJtMDjdM8mzN6LRyuMbNrisVPEJBPI9zA0B6FUq4o6AnQWeUbnpliFgBH2wsRxUzkyf
38kCNBSYeKpM5VULuHumc2E9rVPo/4Y/vRNWPhiha2mt64GLc0PgmvCPoBNgSh7gcjJ8IRFTmJf7
WwhAdtxGNc6/q/XKwxyKcDAGcXAoh/CSLt1hyfZHgn+lBzO/OXVgDJaifgXiQ7rUl1+3DRDtdm9I
KBsqQZnLDbRcwFkZrlkX6HB3AMJnSJl9PwGZiAySkrOlsowxkna1VzFz6ob2KjgKY1krqK9Dj581
Mkok1xX/tLytOMUc37BrrpxAd9Cxy284WmmUi9zUd0qRUybBXYZxyq94ScDXZOXTVbvr7NfK1/pv
D4BG1bdttgDs5UKwQyIyw6ieDgtyI6gUHJ/I9WO9VlLYXLlYMn79pO+0zaYvE6YIyQY8vnUSd2cP
MMUySqsUukMDtsga9Ew6SoF4EB14a79XSLxb1Pj0l9XxyZO0UKWxX0nnHiuGQNY1uw59vchfrGYH
21i9y8XxTaJcu33Y0aWLq5ynYMVx7eZ3c4DJfBJl+6LJ9KNCKsWudYTeBBbhMeQ8gSJOEDuogE1O
VMJ6cMySlUFp7u1DJE9v7I3Gs8EiUKJLMH0kUimEqRF84W3pYZPEPpM+QZ6YfKzl00XBj3lLhE/6
VyA48xCQhKLoqSm+m6ys558jFpud4M4PH7jor/5R7iSNa+9IlnHP3dNJWjboLH1n8lDEe79MmnXE
x2/43unlka+hKBbP3exgZVHbZeSNXqJXnYp90+m95WKZZjj+xDFfdFgOtEtm0Cu3RwxvDA2ymy94
LdcCJVEGf5M4N4natXREULstpROFrLW25AlqHzC6xUTU4QTUEa0XPHQG6nmZWXKwNoduobZUJNGd
OXsdVPcb17/hl6Y7N0qYD55hTqn5bKKppm+n7LdanfcYbGXRS/1B0O70BT19ll1PrrLozmm+/w39
B2pAbh5cdUQfxOigpDGgQMxjgfoOBeVwjgPJ7R4AB3h/4wDwn6kcPpFn6SZGYV7mb+iloXeZhDxW
pKdVNgEVrYlLHi3YwLD7iAn/pFeZSUaqa/k1vWKZ8BrFuhjlYkYOqgLLR3C1ZaeEIU0t256C3Px/
DNvLBjbqj1IwjfcPa8SFWJXUv9bHyG29ShOiXem5j9gzRwMFblWm0GpG7UNPxk6+lBcuv1TC4dYj
ZR8aVVbzAOUp4S81pxll3Y/OJ6kVLUnMxpD8T1WSyjKWlgahdrhufMz8Eu/Rbju1KuBdJOQbLlPo
MVODR0TeivSD6qhCoYVBheTYZ/R2GOi5vm/MaPO5uO74kFINBgUu74yzk34b5r74eDfX76MKZgTK
HLnSAY/OBGvvcTinjPZ5+A5okz6u+t3xbQROGRvN0LezsSn3TbDGXWvtBX+ixCMlH6EZQX7je6+z
NJ2zENzS7RuJJBmUbqTE2AgsVif7GdTfGD3Csis5dCdyVoC7GOt0eZMB8/EAuI0Vi+UCv7B7P71r
xTqa5CLiionQJJNJWo3XggOAOEyaeyegEg9quww4uScZmCKLCl6vcbldRAzQd793HAQYux0s6dIL
NAzcfudEsxXZhSyGXYasfY8JxdZYrVur9+upY5CBCF6AGRHHi62FfGtHbffjm5L83ZZpreGZCMDX
l8UPX0hfiQC+DMjlMxH5aSVGERP2pHaYVTdIogQyLYGQqveNmVbwZIMo0XEA+yR8ORM136U3XqXl
LPcXIVYMRt7zdN/sDi1hckzHaRk6R+Qbe8fx21ZA3xiqoZkuiliFRDQdre+vZrFSkt0bO3TdUTJ7
MnehhClRGw+wEDMgPFJrOxzzyU+7eofYUX/FIzODwC5PG+GwyHxrtdJoVD8T89NWuehdk9AOxfQD
ImvtXuxoC0U/YTJJTwHtxL0pc9qlf1n7xk0xXlDowot8DwQrw9i+mnckwjvxNpwK0GBP8XboCHUO
fDlTo9kfLCNSXYx9z+NASi7m8Nb8f5d6DBRpVDYeqKMQ1VNyGh7ExN6W/7ENkSvefoAA/ysZkH5c
TiFRcoZ7Jch7N0ucL4VfZkWWX+OJjqo23szd1jtQ3DJRdO7PmeiRvwP0rQSlvhdHSsXzWwkX/ACC
DlD/sh0HNzH8Ukem+Yb1C0cY50ukT7xi0AEtxcGE9eszVaBuW8cIC4Ib5HUURAOLCIjvZ4ikjsOb
kVfcAQnyRog2d/8pBLNYRNGw7zB/MmIcsBuvWoda/QFXDABdPxIRwnF0R0+Op0afpXvfXhg6KGyk
ayMrrTq/Kwv3lxvKYlQ09PlBB1VJ9326JYSq1cODcbVZQ3wAmhdW2tYhYTEE0ZDbCRl7Ay6++oLc
jnfUO9ERcYTfY5eCVSGGQawYLJkVZ5V0Q/0jWeFtuCa2rxF+kBYEUdnYa4vW19x99ktGJAd+i3GD
2HvamWmpMPFc4lOvbG0jhRZ6Ai6r/3UzUKceY+FkAqkPv0yTaRTvLxYCEA5j+Kly+grqcOBQbJtz
sZ8nm6wbNUsp7PM5qWMHCQ3ETbJK07Lo8fi9enZf/eKo0kpo+9u34hHItB8DWQ7G//+DBvwPoepq
GnOFO43ZtBsGye8NfEsCV3HevzdHkqDFwZogNJTySXcwumppIWI9m5yL4KU22/O80u5/PWpJmnSk
SoFqXMDSLlZLCCsY8gAMnfzrghojIyIjEVWWPtu47r/6q32+8NPwlbLm3PRDBIltOFHKHG3ZGlc4
38B9jYG5U/MkHPsagz00IleWrsq56clA+SCkGrVfaRa3Gxv76dbQAJdlGtO/bktcLHvLVKohESzq
MJDF5DIfStDYbFwEhduTwycb3GpxlGbUQtcYK+FLJstLEbIUGEPub1Vyb/O7Rqw5ML5WKB7lyYAu
/tC5AqcDByhSne864vRxKXPVhj3fUAjaS9gwnJtrnzCSrPINiNcLVFQxOkyK1W0GvGxZUTDKfhuw
dVfrljAwZgmLtuguQ5V3DraJciG8Ye9qMmeIDHc/6Acv0esXIbQ1pLUxnPTjWZGCmAoJFbsofpFS
9vMQaOQwiy4OdzZ27ilnS1JbLOZdwwoGE1Yqpuml9Wi7Sn6S+AvEeHEd3cV3pJGQoc4fx/eiB3DA
5HcLBSZFyV53OEK1w2O97Q2/jyLUU48d78tTU9ejQ2U8G/BN55QMaVzscT6d4Xvprt9yL6qwdZCy
s+Om4+yFH3mjCtFumLcvgAcR3V8pjFJEsm0MbfUDhQf6U8ZjXgpx5pP8tTxgnNdJNlzMMmXu6tZB
k2RrYq05qpATJoNzGK+DrqwwzcRU6+D3FzvkAwr3iXA547W24brtdjk1EVQLZPiybIF113cDZijL
WKwousO1w0ZWWjRIkgmQvKjBMB4d0tNdCbjeriXpRkEiygNCvcHRlg8NY5/cWW5I6VswricX/O3/
mopEPUM6+ntAFFXlUeCQu5VFcO77RaQPCDeSdBj218Z+KyV5RulTKWmGPqcpTZ69HCJ2J5U7LWAq
WPKtvu610ntnNDc+2TKJVwM6VPNXxGHohkh2hJCVjnKQ9UpVfUwEL1Vp2cqVeDpWQ1+x1+uHeY0j
QXkI+mloTBj3TILjJbtAW8m7BmrYYSrkK+uLE15PG6d0kYikKLUGn21vhvIoB5yYA3fssH0yeOEl
xIJWAEzg9yOUMl0iDK8/dHVmrp/ufukFZesQ94/JFikRC8uvsuIPDuaLbkuJrgJYIQBGpMQkD3tR
5Tz2EuHvh1jC54Uc5vPQbxi2esmnEh6j4UxYkGr7BpCsmVT+N21H4fe0x6LfL6+YMW/HpFWAnuv8
A3kY4rMEhAoInAuQvjPlmihY1iu2j8rJGR8sK1Y+8+UXkQRkSv7zzKxBwfcKPgrVvSLsHQt3/qdv
bReP1b+5ZfoK8xi3wvHyZZgVS8t1Ei7xa3V0b68LtF2tPYwUGnKEZbn0PfZ23oKirc37jGoc0P7K
oYK571maXVHddjOmHE8nHF9XhXmLd9S3V5GpQL9eyn6tqH3Jur7IHB2T7clw9Yn+9T15ebNUZXlB
SeGCEgMKBS3h/rgMiZZsMBaiza9So9zC9JmyhMyyzz0vXMfbGN4ouZrvj+EF6Tn2Ku4Epp74zHMT
GWuEjde9CvNjJPT6EJf+9fhwxexZnXNA6ERlQDvI/57ZenQ93HVaCFgZ1rqzMRO1qnYmCfk6g8W4
F6HNQuiF3C78/RiFFZ/vBmJ2DxnAf3GRUmwyUtjO+HF4CCLjv3+aD6xMq75YUfAdT6IvwgkAsNQW
QAPWwaEQDbCVrkMkO1/qBqdR9P8qQM8hFWfAdGrYBpy8vpcnMI9574huhL0a47XzB+2OxXX92bxN
Gw8MezAq1Kv6j7Er/PPIOlIEE3YW+jpbDkxiDwVxwA5/j4g6Kv3Js7LAmA+p2fTl17fTiYBtsGRd
ofpFgzpVhpwxjW76Gex1IB8gSzM5BeWXE+RTasiZDrgHtiZQKmN7Uldx2DIUwe5c6xas18+NvZv0
aJiYT5yO0i4hoDej+pLABKAGXIM7zz2OCjjZjF3dOAyb7AS8nJEshT98OShx/6ru9+dTx/ftfCYI
kpvcUVDFO5JP1kzlDnEGVQThJY6uH06aH1knr5mfMu4EjNYuCrZEtki5jpGP+CY05ekjjQbNXUYa
ljgt0qlwcEkvz1oRRyINRK0XfVzQsh11KezX5sMWosOxaU0IB/14ZH/28xPUiTXDWd23wGj2PH/A
FPe2a2ZZsM7MB/LSS7GR3g39WAWWTKxqAFA6uam3j0nxQZxPKi/vr5lJkeoyc+BQOk3769IOShsU
boJXekW0hsUH3XjpCk/4XAyANGZMz+7t63JvGDVLZZLVVJkC6c3NMd7A3bKABOEX+Ts1O654rQhi
KyaqjkCXTQMVFWJierHKPnXG/P075WtWJy84EG9vvpORfo8n2fcYIwTcH+W4gyWwSpEMCHe1Us9T
CMNmgCFM2chOzuNXu18MKTyDlSH9o3B0aHkRQ9VXx8Gf3Sqc/mHr9O3nUIEhaLPUMFNd0Ov2C1mW
7gMKmD8mEtrJtisAbr9CGprfRMnZ3Cf2ROWS7rAo5cBVgFeBed6iM5huNmpwszBN2gZ/Lxat62a1
UWHMnS566ZW2SIqIXTQX+PFjLq7DER40B6nolr2ajoRdWlyqi0GR3qcxUVFrUYM9608ePjAbqLAG
N+BmJCKEjpLryxWFSbdfyOfnLdd+s19pIFz/MHari8Tw38HhWfbr0+iMzN+cHkzTI3cUrna50BV2
T7PTVz8nCCszbELU5ptkg4PtOiXwzyuw3QAWG+C46+3fIudHs2+BMXssgfS51vERtp1Rw+YVRYs3
/VVAv4E5ImRuSvqzo3fK0u8gJGcRCxe2h1CJeJMU27r9mueTiF4f1n2MwjEvVDAw9ARHtqnTLDzL
F5FnwD9p1gNvPWB6yFjbzOykQD9qy9WkCwMc6hiheF742+MZl1piyL3dJecl8l6RIB00mSX+a/gU
6yz9jNE7oQ3AhAV3AdzlkeKSTPwDEEnOGejoxJKWVscwOziQCit5J/xhoQmRjPncriyA84DcSrco
c46+teBaR2Dn8PJ5rIfYvE/BM4+iw9PR+Y0IY6n7C9a3njREXffZ89B7RNVOuS0xg4BU5UkS/0ax
X8V1hSEXeBIs//VT5d5O+oX5OXhUElwL/++zoR7pZ404xkkNWIRiKLIkVGqz+SeUlXhdVS6ehGU0
H9j/TMjVbvHAEw4QxGj326NWPb5LxwHyLWEPZGI/kePPgn60+pIYFcApZRrUBN7AbTPhrKMax0g3
fyJ3ASHrIJMJp2tqrorYZDYEQ8CEnJuPiuRZrI3G+UdqRdvZj6+SxSSSNpm/dmAEgISnraq7NBTj
yNrQ7lcpXRjBIYu7zBiM2CDwhALiItns+pQHLmPyiPYr6HuU2aFYU1uSxbTQ1TP1IO8Jicbqu4OU
GtW9huG374SwEZqskDXQLos3W3wYpJH63TTEjOWBSglARIn4aftcPtOFKw7U6lDz8+r2UiumyMKL
rTyPpaV4TBWZL0VIGNVQpP0DfE3GtO0NUDJN7qlAUJ7EhjcY9Yamsct7puj9oPalHv+t+MLvILAA
JKDal/doY6GYfLFFunZeTdwlsMRn9vrGH3vqJW7d9AtrpLailMv89KiaFRpdCKnu548aF7WlI7ST
+RJSe/1WCp8T0XIBeZFtkhL3JIMpf1n1buCFcQoTNQpUPLSwZR0Q2v9/ecldRjA78daLCyC/yOki
ZuQHlE+UILmi/ijkajcr4IBgeQ7j2aL0/FWQNZ4cHxvEtNWOtAdqeOKAOUxsisEz4yMhVpm1UVFI
8LT7Yw+CKbdsRRs5LKP7g1H8k9XCxIe4pWSUg7i/KygIffAT+9mAAZdJpz9iduq9JjFIn1F1jHtU
03wXLz6Jh5mW7oy9SUQetIf7t0NOfkXsOAbrIggpWC5XYTRmT79+Eg/QvGtMFc/+SqGFNhZprjSj
R32NtMwbV91NnJgxdJ0r/E3i6GqoInu+AlMXqeCo0iGW1Muw6T/NTA2tU/yg8CqtHVZTXXqXAzqa
/AUcRRUygODWc0Vb4wbg40QyfhC9O8ZXcigD1K4JBN7fOPn0wx9QSP8p9RldWg1KrieKgi9ks3cx
250yBXsvCDUPze6ZvicY5AJ+trPpf8sjn/WGOJrW24E+t2LyDL81tG1QF6dXBeuRmUe3TumMpUP5
jL/3BvFTC1hmU9nI/qbjsOfr+X9niHC7FuXHay65lLwUGw1gs4MkOGyqUW3PsohuiTIzeBjG+he2
FuBwZzfEdQX9SA/lVWUMnqw+5o3HgLQTNFjHJfTIp7WQniPI2+UjnmWrCYOWzfaIvrfr4D70C7l+
bPzDQBeWdTMHx8NZZ68SIA1xedTZl2bzrdyKm96hucnG8tz8QZb1qCjL+XXtbd7xxAt0ZnjafIWc
sMeFaHEvtfe4YytOTov0475LnP6UKNqJGgLDvSTXobd+OrRF7t2hS3AHoTlLEg0VaLpck8lUaZqk
+8iwnaZc/4XzlZ+xh0Be7bqRWnUXf50XXeDyoBnnsGn0W9SCq5JE413RK05i/kk1UvWvSUqId13W
Qz92f29fXtlcWKoi/fPtiZmh0ROuI4tADtxASDSjHeJW5Hs0UQlhh0VtDaWk0rAymv8YgNk7Ekw1
z+ref5Qk1vcKinX3gumyvm5N9p32aICyCxcEphAySRbcFwPzn3B2wxomblFLFpKg6UkI8UWC7bb2
ZE3HAuYt9EB/iwlTeCGWfQ4LB7/AsIR8Y67fxaW7hs77FoFyZ2rPX7UPabSKtPivXFXPQDK5PEha
2sUK7y2XgCSVBt4xcPmAmQ4Vm5r7hMaUU0BG46xTrRwaqwou9OhSX045wAntuAybmmoaRiVWwH8f
OwJ5zuj5f+y3BRzqkm2UCMJtZHV8LHTo/b+ZKMDQkETrvwJ2IQvEvMViBlfZZ1SK0FTuXzMGw/Gl
KmN6eQEnusahlWhC3JZcr2bRgFNmpRNUJv7RAHXXDf9hq1McDBcp2jNlt/pIg9Wmg+Eoekv1KbM6
L6ig+mIXTA6qSr9W1l2+S99BsV4u6gjJRZHd/N4gRn44pqTEff5euCO5u63l3+ZRTeiqhPA12St4
jN8JNlBKifdh1gsBfXo9gxJoc2YQn2XnWXG4jQu8BcKFUDG2iIsIHGpE7x76QQqqYt3yZpivrjRA
8KsJ6d8YoJRiqLKpesh4ndiiT3jODKx1vkvdd3BiZJxtlkeGeODFgc5AmQikyKws4rtmCo2fhmSb
sLuvGQ2LMH+q7CCTdJPWGpCkHbMTPp3orUIbgKxg21mqY6k2id+VB5+9ExGgqdV/LQRdc51CloQB
e2oeqdbgxmBXsqmuJX4h3vWBGk2CSH4XU6i40xSB6aOFwpBFrO/Q7SeoFng8Z07ilonNUAdjc5OR
JXvMsIzJnk7IrMSoz3BjBOeih5SO7kp50qeSSAd3skgwhUC1I4ohsenjOrGZ8o0eUgj1sdoSHGkH
nYdd8N/jcQ+F77ApslJHVKTQiGnOJt2+DznyL6yDUAxepqGmET/tUoJd2rLcTEoxLzebWm6vs5eJ
V3dsTpb4mAdurWw+kyBR4ifDCK9S0GKTO/2J7753GX/h8OutGH/fR0COQmQH+3n6r1WaFyxnxdeG
xqBZtRgInJ5Cz+snXksh3PwY8kWvtjctRfqWMuj82cuPOFqiSAWVmjKkQnUU/bC4aJh0Y+1bXub1
YlmNkEZQpQhiPT/ae6RcKA+gOSNfnSXQeiKC5h8wuQnHuJdYEcFuWrtqvEfTTkRevPjVzMNWklpa
vaNk8B/XzsUas2+PGlthfqiq4PGBGRhkmLAxYNogB165H//XfPMYudOKHJreNjuqPLEMGwkfXKbn
l8pF/Ovm3otShULw3hESWyU11ujoQ8jNTbyzr56uR9/ZK3d7aa1IKSp48IMdu66Av55mBKh8DkDo
VZ+tqAXF1MwcwhAFshRteuACn4842tfMkeeJqiic9dpEL/mdwBG5VNymWgyw0cGKWHFMmlPGgjX4
YDJPHNe/Bz1BCzdF6DwXdUrpiAIdwFfmD9tLu8fMIS5cPsihVbu3BIiI31/zKyPI4ITjo4zdi7or
Emfr2c2wiim902mvmeeBbPN9XAyw3Sn/5sX5gZHXIZJgD509h4xgm0AOzapEEFMkLLuT/CvphphM
NV2CUGS8BzuH+LDNTuuF0WrOGhG5FPgRf2Yl9mJ7CjydKZnv+pD4vS9ewP2h6/Rms5/h+Zuf+2uF
qMca2YWrHk6yBWr2QYMDHed2XEqycjlq0sZileVCERpZlGxKlefucBGmtAOBTeuO8n+RRl8r4VPP
DQqFHJ83n3eIWlsSWVZaG3AIBSxHuicuYPybacyTeHXDFNX40m/8XqTbVhrvx7GF/9Y++GaAnYtV
QkoTbg1Dl0cHOBD3RQeTOidboDMkt72V//C1Ka8gpf2Y2G98vsQv9KAKkKAgXI6TW9MoQrnCHBon
h/jE8JCiAnwb2eZBk1+icaT9S7gsqQGzZKQtiD8N281Dk5e0ruOXBVUpxK5vN/b6yUtRNdmWIFmX
O6jQ0Z1jQJo5XrZ7IrAUgq9aOGj7Jgtm+joCS5ttgXNUjbErjky095EiT2jIVMu5Eb9wLe/mvgG4
lXS7kb1tD32GrBgVtt3i/4ebBharxR2U+IQ/LLqoAgTEOWwbAbI6x4NC1OwVgshDxVaeMX8pU0f7
CCZz7NyS3WhI+wUh0nkTJQ7E9Khe2+Wr5srlQS1K9mhihH4PvMCj7hDObZqLmBYd6Ks9f6i3hpXw
tzHTGdTCVseJDCweR/+vdf83f5b2y5zvtQ6d/uuAG0wsngLt15ILaTI4ufAfLoOYGr+3RPP+qWRX
PMTz10EMC3ob1nvt356IpUgcNp2sQkxome9Tcu6GnoB8eUiMTtJ5DllPNGYpMZCdzID17/vg7hAi
FmjX7utoe2Nijp99gijfxnX/G4CXOaJuS8J5/PChh+Ub8h4F+HPklv9bAdRNcddlWeKAlGXVCht1
pmmTMkmTjdWhh6ZMCnjP323Oj2MPiOo2KtbpYT6Y6mgG+U2IJ7+kFhMuUWsy62IpV58ZM0oYomM1
fR87UGUMxy7uYwbh/AeVRbczQa++S7Chcm7lUDEBdoALJIeHxDgQKNL/j5mELm6P5GYERC4/iqY/
K7cTAJd35AgmSXOXxvl0+2LMh4g3pGOzxPzLbxaLt3X3ccZbEV/3k3wGqsFqclEgVJoRR8SzdxQf
RX9YjZcbAq5H/OoPgDfb+x7Wv4SEBbpFZpxabeYJgqaPxPFQCdpuNNYBT9KTqS0RUlnmmgVPUcg8
EDryLWdlbyGRmtwPEPSSGnltQruJVGZzlUtMKqo7GOqQysHvqTeM2bKEeZHVZiM6cPXvVcaO9Hj/
GY/iSBWlqlJwUxWaQ+MUre8f08cm5wSFUmkDpR1EGIkVmP96dymeFpmxurtd7JscfSnV8IJ1ZuDm
/3ZAynNXKB8n+ToFToYXvCSANbYWNqI55xEgqyTVj4vH1BaGho0ENWojIY6oG3NmYgdr8vrwbJ6w
dDq6/piEHRTien+75M110Y6z2ObH2hkDFPuzvGrHFZF766mGu9ErDXQc4tl/tUaimg0Sk1ERnZwi
0uGSjATCCzq8Q7sGVrKCtxfjaZyjG0QngOcikfKQhDS6tGfdAqD1sAMTisiPIMClPnpnJk3k5jb+
tu9DJ74yfV8YFdy+uw+9C1dIyzzEe64Kn2sUlSgpaz5ytq6GZZ/Cegsye2uFSCG5Hb2puDIdRkD7
wGre5M0oU38NF84p9xoGhIgeiIF59GR78nznbv628mkgVsDQFa19ShaJEF1IFXmf2n9/CWgnTw1D
Y6/A7f8P+yuk9oIKHqEIGmQ2EFcdGFm0Iz3itrGQC0lDQswHIpZXLAc2n+L4RXBLoyiHvBigHLHp
HPRsBi1ZsjYabXPdAM27sMwnWEUNJF6VZxN0yN1HZpOfgTa+ucvgVARA8oyBt07PiIwkK/YQilyh
6kdqSQjfDgsROS4+6Werl6a5eu3pLs9ko3+0pBhkchHmMIJrIMv9B2rlRvU8rT6/QGHsgMDaO55B
VkIJwdmIVg7o/Mp6btqI4DpedLlinx3IJd0ng3Cym9pA2ExPGUMhn07puIGZ17YZSb/l4d7ANf/7
doUD2OGZHpjm7LjGwznAyu4EqTM/Uv456pZr2MncIMg3PFhoHN+7k0cWd1RTiSO/TVYlfpQ2FgIX
S4PVpYomVieM7pOAmiMKyt5aEwFpxtdd6T79nN/bFtD6OOMoBxDUOdCTnMdJeCfvmOycwZ3KZO8Q
/lSPqY8zzzf/9BAOdvjo6SSKfEEx4Kgl5TRYeSP83yQN5DTG/3GclLRX/SJYUJ4SwJTbfakD1Pfz
zezkc6xL0b3dXBaYBqIxIzJKbvLcVJa1XmmS9XW+h+e7Yum8G5Xy2EGjzmKdeQV1Eua0KZ431NzG
vsF66e4qDEYmiXnyjbPfIkzSoQuqpvTbJZXnfzryYKoIvfIYHagHo3xm2zD4D6LZbY/5x/GJvMx7
GC/sKXsdT7tYYGxt3RcZamf8J797839L7EAXSOlFV/raw3V6zlPCiEI20TyhzOg0pK8+Zz9NxNTH
LxiYWw3v8sLGgYUCTdQdSQB8np/GH8WmhvXI2blyEFjWjqHy/yx63WavFAlkdY+MwaLjbvKXsUfZ
p5NogDWF78YZVkNa9Basf+w7CPqD5mYIj10uHq5NwcMjj3tQTAqJi+CjNd0EJl6E8k+p5js283mu
MMElN6g6t11qIZvk5neaKZH2R66EF7vrtIAbj2VWcM24lbolz5I9EQJxBEvlYauh9FHL+BGpQS58
eXcv4/AUuu0FqKXiumWX7Z3Bfbq80icRNad6WNmCZHPX3c2uf9Fj1neZC+nLF01mzrTB8b0J3L5g
FXSu2P/9NuLjZrp/T9j5ACFLbyvUdIfzvhUtnofWhlCMsWuth3Y2RzG7QJQMqppA8jvUDrUKTUKs
5CXbIn2FEGDlJG4mvJlg81vUdLzTBUxazuALPP5pWJ86Nc792dSN6LtZbyB9B16fOgxdQhCGzxty
XDH5/tpxItBel+AN14SUUCopPMi3pep/tAcreuO39NTtVqw7Vsw+5/fusvynTby8e0Js/cPwdNFT
5JiHHEsdkzsmFDTAXnbRkJ/maz+mWTaMKVTw4QYZCPUcPQXPf/cYp2Npm/6kXlTKAGOX6rEw28QC
hKKsztUbYKkBW0BgQ0jNBdwqgQXIdomay5Sw9UJa+eom9TpxHr1ZccuWZlIQuFbeFdXhnxWAC79y
V0uDGWKteB+rfAeFKrpwwffYr7m3K7e6zAYuqKwSb4yz3hFZnreamqVb2dxJzQ0hI38JUdSVx6Sr
etkAgDYUrUlMykdkaoi2GXAOr+oRsT6FlZWEvpsmNNCVCIZUy4OXp+vwG01eguAa9oZGHIW1JXzS
gDaDB8eehn85ElqmH77WdIC6ALWKMrzonfGqgG1i2aiMX54IRFEmu9X9DEvUND8jWcTRoecvyZra
WER/dGMRw2mklLvoatD66qQnocyNCln+M6IDv3qhgeZmZdtc1JfggReOKKpItreZ9GYI2VW73WLA
H5b/sWIVmicEnAonPJCy7YC1u2beUNixUQ/oteaN4o+Dlq8UyDA/VbQEwCpDvWAY+v95zEym1lN6
hLZtrXatsYI1z0f+5rdkFXvgJuHTghHR8XDP2J7h1O6SDeOOrmSjKkPtD2VOYTK84Sd5aO8vdNAk
tMRTA8RFIpHJedWyvuzCmlenHDfFfyB36nyDNRCEMUMZgYm+ur3xVVheBWU7I8PLT8DXe5xeISbx
5jkqTlMOjY1nnGQ6h+3je2Cfdx8UvlRVL3akJcnuVSoJtLXzA14nNmxDZF0SIpUja5q2cB9Uulvl
u4yHFahLaFQDAz8IffkoPdpUb9aDlVoySgqTYLtrdZNYlcwvUvx0z5IWgJEoLGVEaOzTU2M3rFH/
MJmh9tuWQZs9Fw16hGSrjMHzPvkpNNsXTRFK4F+F1YXKWzmcMUDY9YM3EHwTJBJ4w+ozvgXqg1o5
E/wXWhL6y22tm0nkrOSOMZYt9Tqcmxg3hdl0nSDJc4q2rh4cbTYyBXPyd/3RMM/UfccsTWTfgYv9
TW/omDprRG1hZuepJHk15RR+AlrF26g8tMGhoW6afXeMaSV1QPS6nFgDoG47U6ruupbksQwJUgXE
vkEsT3agk282H6I7EN7Z+fgfbcPDMh3VfJWRWnihiHjXOrx5FUFp26++NErg5S58z9mc/scQOGhV
0x12qnDYtjLOWZwBMUoWShh9Tkj7sYrKubPNg9e49LhWsuIvPfSY94OiZft3Q4wBkCh/XSWa37kN
+zwOi7Eu1yNwwJINGnPn4aKW6tCJI0R65FMB01nPZIXXh3UJMUdcwghDCwI9rrrc9zdysu6fTn2l
lEYfQuDNE5dz/2JGezI517XqoskzsRKMLffWVBY+IZ1+lsj9HzOEbkV6DvtSr1yTmSrfNjpTd9ca
+O7Y6w87gsOYaHYUiSTz0ETEY6TnBNG1cr2U5/hRDCYMrn1xVe/xlhD/6ArZx50tyJWRYpoUKynA
YEyFd8i61FOgbcq1YAFsG0PyCXQWgKRO59bE3IOBmy0ndlY8b4KTYipqAeGUHiIW+TNuGFMNp0YO
uS1SYjUUtz5DzKdzvaS+3aWurzu9VmqO7dp2ijkM7KRGT75hE5K6lWlxxpQXikZMK2Dgh/j4d6pO
AO70gEvvS+GvAeF1R0HtPuBU7bHoUjuBH17CTmAzGp2f8T0rcPYm28qaAQcXFkgGMyX5Ss2Ssyvy
+UMHCKIMGQMSZa3l1pQzeHBWbMHzlvEfsycTw1TcIrtOcidAJumtCFUmIYBhYZ0dgUxxBqExpRhR
M4Cn4vbFcUNmEeBju00xRTMXPPQqShnhdHJyOtDC2jJEP7tFBSl/83z2HYTR+G7sZdsSYmiQv1Kr
/9dcD1JWi9EW2XkHOLXzu4PolgiiD8HutGhDYPG4M6n5qLdFXRfqkXy7nqstLAKGD/wnmxUV9bdj
qHQmLsxZeqVNIgR8015v896sZmDHaG6Iwck0ysvnD74Xfn37u6JPX+uKktbW57sionT3wriTQ0wX
06ZzS+He3pYWfeAbI3JR2eBomkSpr5K/JmQ4OEwdrBeEANpOnxw9YuCGmBAvu57vsAvl7h2t+lgW
nDKAjbPf6KZ5dmd5Vae6151asI96jfGmypGgPytuysbpCj8Yhng9GzR4XW/3T0laW3HY+vOdARPB
BdwE8x/hsM1Mv9MS5f4SrkAwsA7FkJlBIs8zhq1o5byUnyCNIOmAalwWOxnmoLxkYUd5Ax4XgMHd
CrggPuX4OQ97nrn1j+d/uYZtuBkkciWY5N8V+nhNR6z6+4D6T1ryUIWgFb+BFroB6So8GgycCkzg
PRSlzU7IExNFdV7BQi1MklgbFL2NuYHjWaFwS+SHjC6XM9xwBjTxJqnZMkGEC6UNgQHDVM3SZ39U
SfOgoDdg22npaPWZdsh3RvyTs4ZCh6kEHUv5C6Gk1aCTBqz7pr2xsIXHmVg1VOcTx5npXIC7I3Ow
TaTCQsjloa2fBIwHb17xJj7Ka10AZ0TRaZxzFndqhITuy2H00JjQXTug4e8Og5WmtIMhItec48XZ
KWP3UPY4JH6E9um5c3oqGKgAeTUEREmcXSfKuLL6k4QdtoyOnF/s4g7LM6M9A2BJvN4OQglvsetX
68MOZ0CbARcfzWu0WMMnitw4qNqVhWvZzlIHpHwDhSyUqrOgbbL57Q8U2yplQ5lswM30G9Bz/5cH
RgO/0eHH7lzWxb7ptsr7TgEnDeJWNNToWGJFEplZeGjQVwGjWGVMmLCzKf36ezxzpRdcveTR1hiA
DBF3wKBTLUNqy40Wt9He17MrXDoibfahICt4bTDQ44I08VBaq/Ub73wydZna+ztgJ6zNU673i/S2
8dWQIBP+HFhsoMdtNULg7bUrtcUFtGREm9LxOlbhHObR8M79aPPRTAynOxHXUFGYWApUR+b5erCf
PmtPC8SnJ9og2ndUXsXV3tBq3jfWOevjpCXHHQANYv9jRcJ6GYta+z7BB2L9tx4XLivkZguJ80GO
5wmkwn0R+QoinH4kA9HpBoNw0Y9URvNcX5L9wEoa5dL/gMU53wdJNumvLGb+eDWK4lr/o7/DgJiL
b0JyuDECvXYNjPJVm2sjE8dYOUjqTVRlkKcaCURRB4xisgm3iJKpJseuMYccY5CIkYqWVk+SARR4
1x1E6M/UGPI292wP9uYk61IaWkdhA7XMGvl7URc3Xbpfiw+O3bmfzLvns/ERY5ORWBBkIFEo/05V
6ETVQE+MH8f1/dQqQYaOi1qPQ4FIfCpnTLk9uIn47bn9Gig4YBMTvalaum2kgEXbYS0y2dHNQSBb
qVIJ1TfcVj/X+5w8ngmpFzh7JL9tLd4P2AJo9TcCwaeUwI3b17IMFSwyfMzla4hshpjvP/3XaLoe
WcBKtXjpu659FIJNyOS147j+rpx60puFM9f4+EgAl3I/0dt33CqAma2yVXJ+9epuyr222kU1ozqY
yob4cLHQhO78j25rLyJ3yeb79piAsRTgc98GBJQNsbSBmrMebVHsP8n0y59/WE5XKcsRHNHNkNd5
p85aeWU5FZ+4SAIlcCFogkbKbmHHtZSmz6L5t6F0rHtTdJdYuEr/Tt8QZdoV9WYJ9zhGorKWLult
SEwWQnOklzZzJkkZsCvv+G3S1q3Xb7kPlBXVwgLrNNrv8JEQtfnFl/AldZBx8EVAYwho1i2LcLID
HeDV5xyCGdcpPO8I+hcNuSSsFYY96471VILOI1BcLYvmD+yHKEqk2Y2MZ5sa+qPNNc1rxzyHQz+N
9aTe5/2CiWOtnoa4xebP9ThkDHqWWIY71N79wmVId2iQJLhEDU8GV4u8vN2hIzlxJ9JCtUSu451N
XlFddWHTH4hnERS2lb4ah/i43og881ZoOiLRUb1GSO4QHwRsT1wUpmvy0BtA8P3a9DQ2PWItH9lk
YeNUVovy6n+HHaouQPWIqSLJEKhVKdtF1WEEuNRij9cw6PD99++pEXFoYTSHqGBpkQJeSYZMP2UV
6cQ8XJVCi6cnGd1jqvDJdOe2VZVRDEorpluP6NxyPGiFiS6uqQciOqCUJyYE0p6la1m3N91uiX7g
+w7mESAN63FOIPsHWkhU4OrfygroWvyJ/LU1DA0iOax5IWi4ji02NDb9WjgejIvSnZuXVMMBDJ9t
R6T9V2FATBt9WgHgvjui+XDQEKQW7eJHGIPv9o+gUyOfWbUPOHVNxll+e3wdvJdS3ftB9NCt/1t9
KYrbL3IpVlC5r95yPTPEE6lWmFmZnxdKkF0ArcmE1iEyD1HmrMo/eDM91hAxguEHGrrh6pKDxy1B
bWAtbgH0GtMzuZYK2oqoO5CghJW96eNTMALiY1npAltsS8Jm5b8pqqzHjez1+XleW4+t1AZrmGvE
F0ocCpeOK/cNJ/lc0G2ALEEasF3TVZJIwGQxyV5xsX9MaPi4dVTZTwJ3RLVbWmYIpM03PURTlnnn
q7NxXv4fm8XP1uMLVg2kQWgd4wAwABqOPmynf8Gk8eJvEsk2qGQXJAdMB5MQbJnRa+GExm1qxk6+
slzW0DXTFwTFgm66v22TGeViverUI4q0K5KFmt9L1H1cY1cAGbKIz6GHlfT688d9fXdxappwmysX
1hA53eEdy+7aVcjSghZ0p8id60tqJNYnGWIIbK9bPkxCzIudhrdMKk87OrsVh5CVbmlHxXWGyOsE
5tDcixZw3tI+9ApC0Bz9zp4YmtWIBQa5R9cviJv+EUS25pZV82zc+brFADZz5w7U/TCE5OrP4QZg
6oUkxeDepUg5RpTaVAbMV5v4KUiicMbZR/zIlr/zb4EnP3yqJqQ9lB7vdlQx7NzbZr8S9pZ0cEZZ
MAUh2y1cCroh7zf7TeMRn8Hko/lcX2gUNu18DHGLa8HhC+T2gD2K8Pt3CDJGZ0bfbKBRBliPOPSV
fkQB8AMRYcyc9gfqy7CXJzXbstB9C4SFi7N4J4qKmWji9oyXwkmdl0Yw9A8H/iMZJfYfmr6UokF3
sAafJ6+ERgmnVIPOGhpYQ5Z3MIub8xWLPFzzWTiMyXOm7KQ04UePR5Vsg2DNJXFYWE12alIXUi4S
Tc06ganQOr/g7T2Cy0Usa8SGTzu32rHvVn3hvvywZvAosdUmGcTYYh6OKbdw395L0plV7tbDfuB7
MvC1E5eJZV+NhqHu2ZPrxUI4M22ZQM6k2iwWg0zxV/UgjLgtM4UIvH+QWkQZ0FLJLXJ6Q9xsxVTV
EbvRaru2L/WCTx3RFhufRPBRVnLzPD/xctth0xt41GO0MEJYG+vfI1NgLCxmobvJrgDW9EvBHmf6
Nn1wfwEIjkbUfAGathpCo/+BOVxIS6DKuUegAKwRjZJvf8ZJALxcM+kIe8EUm4DtCXD5lzPbuVjO
ypliuNe1GowY17T5Kg2pqrYqIO1DWPzcTZFfIkex+fqv8fpJY9x27LI8JVdvnJC8Kpnro99KF1CQ
NR44kVklhZXfFL1FxdoRjhARmOPBPEGo9G/QKx5fInut8VZPRlRTiB1QDnJepMbibvUuVRIbyMH3
sZ14KiouMbTx+Esqhn1JeR9ZgB9dk7aqlD371ZLtDouVQpv6NNwHLj4cLIJTolAfU5ayyf4IiagY
LoIB9nB5FEcrtLLPoetQrlgeuldmGwio4NXdFDaP8UTC/ntaKcLUffhqYr3vUaC+5HoUhA960Yf2
kxDZ49xZaWg0DipGL9UjdkRny+acmmC3lSUNFD1yBurXhsFU8URQMFvtf7c4S0bmsnrXFzA6J1aa
o+HDQsQtUKErR4E3VBO3FQ9Hqg2f53FAMk/cfgcb/84XpcRMLkOXoYi3rukJP8wmYAGTrquQtA40
VkufCSeOphLyS//DBKF1E+scd8VrDcdtYkULhwH3q/cr3K4Nx3QSNXEkAc4MtQICy7Gyq17LbeOs
FI2iapIMqC6RsfdwU+rEDTAF3JObLNv/15W8jPXmcd21T4nVDYYQ4CcQEmvJeya9NGtQkzSMG7xZ
61V/f9gUjCg8pfykCcWrtUk2pHXOAQtEaAIwWfRsX5kYPfR+q85WXpAUtqYvON2X4JLVsFzu7o/+
8AzDYZiSnU8CluH0/MSPQE7Ur7jqIuO0nJIQ4F/Hl4Lh7m9iJer7258PUcZSHmX0Zojx9jO2+XCQ
9xACzynp7Il7rG5qiQF+Nh9wPzrPa7dgkdWODLZ/Bei4LQS5qRlL653iXyI3/qTGWc8OKJeV3rkQ
znKxxfWDvqK78AEuiAbiUym0hTBoiEpqDgIZKyg8aHBmKugejMj830bY585fDI9HKiJVEC3vDZpO
n+6bNlgS8/M/BC9aco60fvbpkfcK1PvsH4cnBJcLkEVfZ8dz12XZKG521tkOWbwCHafF/EdfdILI
x/6Q/8KQQ+lJlyfSQ8iA9qZ17JljmKIyvGhddQlsipWRm7wJrw6R6TMDj4dFIrwdLbp6cTBp6KzH
aFNs+IVWU0AnnKBK+OE37mgXAPTnn6Hdteu2Q7/OMmPFWjjuC5BMInp3PYop1u7PxN3qkbqL1749
td0LgnmbLlc1n8DJQ+FV7o/p1EOiBfoWbLJXsMtjz952FT5X682ari6JiDUmGHhUzSUXtKqWDNXF
4mJxIZqco9B+JzJlxPdCFuyiYpam/DMxeu9fjUVcOY6uROU4z/MWPqc9UjcLgBZEZC63HfD0DeCi
PGJGremiSZc+za8Pvsw2sTcWg328pNibpXAYrbNOIf/HxNCi2plz5y8ltfFoKwSPH0hP/1cT9uod
2ueIzMD2eAkDkWI1UpYbKRLmmUFmTWyrVcd3oL4T9T195WH8s8N77KkCuYoZJAVf9rl7qOEvtbFU
2hqBEFioDifTEt/4xmDzhot+BMI9Vz5c7E4IIfEodWd7rxbDEP5B04YSrYugEY9yRo8lS6c4/uYn
lmXBxIfE1dd1szrbF6TAfWyQ2slo6lh8IWF67Ex+KCOV5jY/PrbqT66RcnD0yqYfmdlC9vbgxCmn
nDj148O38cX30lgvl7gfKN3De4yJQHD+Azz8u0BX43jG3/65dfAadJ6LMaiM5GvYI22Z75QIdNXD
vY4LCgpbCW7ZqkWSw6rFjw+pIsYK823xbJ31N3z+xe/7UeMULgLaG2PeSN1JWzIAt96y15kyUwBj
fztxnqlCQWGZVcp10ef7LdBWYGj+dqE4DKh+d2M/dwKul0bKnX6+8nSQ76iozeZiBAFfy63zK0zL
NWSZnofjaYCwu73KhzSkTP19TRZdY3Rq+JOVvFYV0dr989zMiOxwkeWsZH4XP8EFqVNXPwyUq2dP
Py2dvvaWsqrr/Bw4WC7FVGGVCaov8BtGvsZ+mJ9CVcitvdysvIwDdiMd1fWl3NpmtgqT5MjgU/Ss
ud8tfaZJqhx9BpyigDIzBkcKpv6mOappjhClBcpbPiNmRATlDM7fhFqc4/MqKGUiJDS3CmoAo79z
P4B7femb0XZySqv2Q2XyPLB0Pt+ZQQyeRKiCr6LsHmH/w/PGoM9z5YUzAHsG1BsNTsKKgxzWEh9T
lpDiJvwX+x8xPJPLoiobijpEKpU+N0xLJoRhNnZLcCDnyrL5kUXzOE21vtu7xVnMcnLp7ye1Q/GV
8j4//Iwb+Qyq8SiGfDP8YJBpBPoPSaKXeghG/Z20U2gf5eURCkqjs3DO8mxJob7Cyq5xPXzOCqS6
7ozH4ayDJ6dKqtBT/PrUHaMQQmqc05RAS1KovWjMn7SRv0+Czb5PT/16FgB3+TjM0rjuD3RV/8hN
jya4BnT9mrs4VgU2H673ZoZERrRQNPYfzRe4obtjz8/5NqciaKmbIpUNRF3WBfbfPbiGZls9j4Y3
pvs79aTk8pKJLmDXC7nNhx6UJKC/d5Mn4tW15sG49WMrwFxen3MBUw0IhfyLwbT05Eb6aAcINQw1
dOLzn32jKZjBziHf1nbpSMwNf6biV0Z5tisafZutkiXLAa4iOUaHlbN8X6MEnZ2AQdpaZAwyKbG0
7f3etxXiRP+YQ4alLnpGL7mu2rgtqCaQyleGEjOh1qUUp6X1cGOWnWtosO4aa4Jp8OWhs+Z0A41q
8djJ0uZdc/RrdnC9o+iNPZAIEj3MEZoampxCKx3U7gmVi5yXdGo4oIYhu6+nknFpP1LNZVKrPgM2
lH/5noflH64khtyv5Qu7lDEgdbL6Jumt0YTo8LzqekilKeHoJqRtDGTMmtK0/cXR6Y/xVn4HQqW4
/tudvyEh7mpho40/ToM7LIWSUs6PtsMYXgBnce3rGhEEXDrLD1fkQBxyYG0a4Hszm/i+zGWVL5V9
imJkxAy88UumFa0K7OrD+nI3U00Z/z1fJIBzXFUlNByBEEB77K3m/q+KeI+uT5LKvH4UPNSngyxL
88KT1yqKpmF2CvOzcDAyKx5y9i3IFME/hg9ChH+jS/hyE8FJgFaRZ7VsD/3OGvDB9TWpzQ79KzWN
Q7dDPUmIi5Y/NGvhJfyKh+v0AV5SrxSwf40mXCN3W8nN5zG3w7bM6NiMELJdDq3vkk3UBe8SO4jK
O7HEj2XODLm/I8SBPPwdfv2G11hN/H7k+jrtjr69bte7vUsbhxT1ofg8iGU7gd5v6+0b86R1AmJw
AvUBXeu86x/Ovsvg9+skBmV/YkY1uHI9z27oeGXt5muCrzt/izM9KY21Q0I9g7Fg47iakq9p4pBP
eNrRkN09FdUqJmY9yxy7DAKmaumuwUkj5TXXd6oatR4cZBb3bXeIchaFeDyqaJMbC6kJljh9nCUN
yM0VQELTbIHi3/YdnWHXqb7XwbZEaSgQEZTyRUeBjBteReTemcIKdgkpJMRrMZZ/7v6gSIVii40p
lY889MHOp4lF5eFX7KA9sVITiZ7yA7JGP+m+Li9ZE7z+jrQJ+vOYtsEZ3yH8GKUQU2I8HdlK4E2e
DXJqVrMXa5RT400F++S5pSnqRo0+KE/NgWZ6rTKGOMRKERRWevjUWMYdCdUOdUw7+54tYvfEo8ml
VB/n33zBWFGc/5QooxTtcXJ98AvglFcl2ytW1SJGmejS/OnB8GL3b1K0madd+osPOP4vReNGQS4X
RJNfzqM9VOcRFWHH8TyalkhYZrsb361ImFlnqYEWG4lRJ7hVDlprIFBioQZCkie9ZYjP1psCJYnF
Ljscez9NEowlka9tv0S1rz7O1MCN/AGqR6N7OSXTBgXitTlEltuTm6I3qym7DlWQknOmz2qOk/iM
sr69fpYCn+ylbh0K+J9xaKaFDUvdEeaaLckDJeB0qV6iugTCrtZOF0MMs73GDAANCJMLeVtsQddB
NBVzkQBvl7lhBEtQ+53bDfO7AKjy0OLUMp9jw/cyXCXXK6C5L8qH8DDYLET5Obuh1poB8YD7Hghu
wMXOoAUjZN/PWLNpgva7XMUgBzNaI0v+YKx3JbB1dJ965lwLTuFkJYgV5IFB2+9UWUrn+sPd7U+w
yqePx2PQ6gV74O4G7PfORKDVkRfYEW327Pyh7aph8ZWDTSQT/7nok1aL0In2jncVUqsvbvVskChq
1hFY2sC4Gtnb8ZfjVm+X2wV4yD6l3zp/RKLtfZMLcKGytGHjK+FC/ytEWsf3BGb+NdjBC2lGm0ag
mDwhF5jnVn/QEo6dUj4IG4x7EiW5ffzj00O97pIvMw7MzYo3QP67AU90+ivh/5rQXu7bkncSSNAz
c6yxikJynWaCHnQR354DZ6aYgY/sxsVmFHYSDoGOzHMj46V9pZ3b3SAxej3SPsZg/WSRThdUTZTP
7qjjLTK3jb7NLp4Rbh6Qff2rRE1RnYFCAirhzkFgxL0xfAw/sRK2hnMenv075lRlCSgAw/vxoSiX
Y6Hdzn58WU8YM0Q/kCKAdK7yGLjoDJMZ0X4u258sOgK2RcNwZNh2OPb93ExwXa0vI4ineoZog+TW
l3+B/yc+oht0BsyjunQihEPzFJSkbpdm99NhGg5kMFH/vL56eIFdzLZTB6niCJZyvA4SS33UhUxF
/pcaX7/qOlXhPIDO8b9DFkk8/9t4HrQvhESw6EEx5R6HuFkMkMm9HO4lxo8O0YLxmugbH1FT1vx+
cSCt0ts30Rz8HSF2d2X5TakbCSsBaEJ+8eFWeh46pE4MBSyQwgrWqj/SEUVZYBXhJnFXyKHjJN2k
+C52hrjrDvwWUsupjB5v2H0HKU02KizCsuOF/ykjAuWfBC0ZU1aykwr0plcnYVZF++sAEhFEb8ze
+8aueO6PophclLXBgZQktirSWozDUJB7T/2OaH+RFk6kECVNyc1Por24BsaA1EybtJBx+0vZHfzP
Hh2iYNLUnyfCOVMXD6njZQqlylYuuY5howiNVPyrc5Dc3+hhow3YswVViNas5GAuVsfykmGe7GwO
xkACSt0iNa79MxuEyLWx5geLU9Kc1wIDkHr6H1NZe5Y9EI7R2d4r6hE39rSWGWLimyO37BqOdT72
QKBe2i8JmDCcOeBOqg4SfjxoNPFS/E616rD9t3TnYDdzUZMqib7IrnV2ATGKfAvnmtjCr6m2GIbU
wTLOJP5bIjTZxx9J3YHgEBuyofBIXOlFxr9Uxv3JQt6OqkCi6FDNVpSettP4YwqCM1j4WIbMuyLq
LdomxL8p60YtdJ3WxE9R9vpY9ra3sHm0M7NNjzE9OoW+NYNI/pSjwzeokZOioEFIxQgpGM2FImPb
l3I7aCZRhtvFEPGIf7Hr8VLL35yiO0Xi0MMZ0QZG2HtDrXCi5ZNWR9QhgdidT6FjxLS69zLxtNoa
g5cZ9gluJqJBWUAdrFl3qYUHM4JDLzrxLnlMoy4OHf2xP+wtz61oJnzwePkhx0fCP88yn8XABi7p
NC73YeCQQ/Q/xLyAusajyQTPoVcdVHhzqFp+5dWdZyAGU9Di2jkZ+p8r6PSuIwQ7xnEdxjfkjuth
VTD7jy7MjQvdcFoQDjmukcQSCeOLBNPxB+DGaz7jtxrD0AaQL6UeqliUpZgomXiEzU/PjgdUMzMJ
aqilFC82OjYRPPfYgF8ohJptfm8LDUy0Kg34pKBXApD0mFYDWlyErdiFpDfWZjfvlgc71gXCkVGa
Vw2eGIDBkqTGzU8wRXn5dkvDs6U1I6fA3CfqUiIYF/jMl8kubU+UwN3ik+tvxkdlw+uOFqmxh4Fg
7qJijHQn2TfE+bv6vLRMLWD5X6gUAeXhRw600hiDMcE8VEuQGPVA1zjjJgqaXdg4PuBBoQzkz7Oj
rt5kO81mgviuBfzhCM9s9Cun+UfKCsPXau2l/0l07LxecXwD83uqnnvzG+imKTO0sDMMqpQV8CVJ
nQ4hU6DMsSGvWq6efFi0ROkbV2fOIzoOI5J78NplPoNj2rqUXJTs/EntthZ7oaSBoPZJ4MmD4AKV
JaSohwzDu6Yd5e4XedRvkvP4g4FWM4yS0tYgZf3BNu6W6ix+82AwyyWmQJvd8tPK1V+QsW6dqKzj
NnIXORW80XpBQQMvUJjmgfZx0AbqoAkzRh15/Je7rzSWU+v6UnKS0y4ohYinG2jV4YpdxF3zGN8f
J4/WTlRN+VFstZ87DQvUdanrBI9ASkDJtB7vMd5C8nd4mPHhakUcxmoB8scnnd+hwCPpnihqTH8T
kkYAJk3WHGeOg+qz0NsdHoyt800yBtX+QXgQ3b8Kj/DhfO/dULIgniq/YujgLtRpuCH6xyQbkH2f
hC0Dv7Qi+jLur6Oqd9lnDdLE/IWiaVWkUi4LG5IvjzZ8u+JkaQ1LoG2/FyRxdjlNbmvSPRtpk4er
0VeG6yLV3OHYBP9Ws1GU6Rvi/GMHIZR07Xe6MJqPvxz/hYBEic5aO5ZJ0vNmEQ1+8TZ+pd2LDEzK
S0j4GWgSqhGVVR5koBqKzmkNHfE7nY19MUH9R8ybft//jpGcG1fydVJK5A6acfaaIa1Fv+w7vz74
SRFxC6iwnGqvE30bcrJlhOrqM4VHK6/3kuGeM2lNV2QoSZ0yQchm6+HLCQ5+WLcBRy+OmhEG/sqf
H2BAwLyBmoW/ViMEOHuHWNwmaCUBJO/txK/DKZGeOeQhWI0pJYyD6g/ew9YU4ol9lKLzi7yq2781
VBL/mRe5VWj2CkOhXj2ZuudzvZdCVViNgTNhAqNKf61rU60TVn0zEzlxTOOyNHG7HwcIYKiVwimf
KnOjEJXejWyNgMzfKAYkizzF35zaVWISLNa0drQsh0BxnBI5RnaL3WSxxq7Tkj5CLa0sV8SQ/5CA
mEg1k7YWuQRg/UhsvFY3a485EijNWBiQTke70CLoXYoLQeH6xuUGmNzQbZfUGTNv8Of0zamWMYv6
7trgkrSrS9Jrsb7Cldg29e6N5YQUHtBW/Jf6PwJzu8D988grtJiPtUZRz/0JdL8q2yzLCh4aOcuQ
vD8kU/ogELPnpDypbJJrHEXukKqSx6ZeWmN3P5C/QIsRojqoMKx0uPV/NFuYg5NEBy49hgiDCNh/
AiXt+HiKbBRd1pEMpqEmGOL3s2MkjmI8QCJZSYzG33J4AuWN+K/TAWaUEQS0rZCGGtq3kkptLQXN
KmPstdRf4FKjQuYorzK+jNnjgx64gUTyE+3w5sFRO4PvEuin/zBuKXXm0ZWn3RC6ncKfGLC4anz6
O6RNc3gEnNblOHTvRgmwwRVPKqIfyVwexBu1858fZeu5n4SEnWaeVZa9QC5zcU8xhDt0O3Cv9bgz
kVC87fPEacLqmM/hBQiOvSo/58GjKr0dIj5To8FtRkF8zMFg6CUZe8TbfTeYyPWH30kq1qHQVhjR
szBKTIxRsTG3VB5QmlttzT4S0F2uCljEbWqRujF/Tdr3QIQW72+wQHh1jqGDnbGJj6ye0SnZscXv
K/wtoHzRk47BHoFIz4ZxyBVY7E+zfaWaqKENn3Ed+z5AxGNMsyUTRT8pHGPSY88w9L90PRTQtChH
npVS+QthOsV/aOBT0RgDnOtvdoQDUGQEWFRgJZ61x6jXHhTrAoKr6Wj9uc+ZOu7NW+zrOGZcxUTx
UVYEB2O9bLod0/Hs5ssbOW+wfxQpbMPFq6J2NLzkXZDrINg9nY5/E2ZFCwLYen/Lwr6tHMVSTk1n
aCze5OQCKyRc5Ihl6d03mOnDPhEB3iQt08z+s3e6xXx9H4VjTYUwE1DVt3lgzehk20I/bRjQCGQ9
yTbN1Nb1LVdpzQk0PPf8NTL/WZN1P7YpYvyOA0HZ8KVQtn5GRB1Gde33mcfAsL1gm9DbY0S9lA74
JE+Ip5MLJ01KShTP9rHL+yxf+v29t8+8mzr5wkz/0MypH2qzSXjvR+ss1NCNHlOSzb6lAQBGe6ki
vXsD7BTftKrqwDRGy/t/Pj4lhPUMyn7g0fr5AerKJ2iwijCUEcMTc6sygE4hugeb3t2JBG1pFdVO
oZkeTFS4os5+q8d3aKflbyVFFPgAPwKvS7tDSN535LyXPAjMLKOVRGpmlZAWpqilJPElN1EeBVg0
BggSaA5ygBwvVew59T9bYGxBEzLZohcJRCwzRJefn1aiVGYff6PTKpn834/uxXXXYzM+egHT1tk6
lMKy3rl92xMouXEPe091RIjGU7zY5wmyfzUVaAxzdOQA2UdVelHm56dxjdxDqYfMp5OMLnW3Kv21
KRsudXS4NXCX4FclQeVMjG/RA7R8gMQzLBkOBVwoy5zIGn8rRGhXSqpdd0jmel51ChSv0H3S7auI
OXzS+L31LhIK/qHBwdWCWnJuoInGOYvSvI8ByWSSmizCGdzkzfmzE8c1WhQAYpVWDePj7ogkRgfT
05zJCZjduqi+oHrlM6IXjG/bic8NyqHm+up+46hu/l8TEpHYCxvR7oT+RMckLpuGvE5HV97EVwX+
13c7fB3UHCsSMm59tQKpOZQljgmClAT7CS/z7WruPZc9tg2EDPaNAddT9+V+NIhDljrPhgt/GFXe
IJEc/Bmv9T3d+/Tx+1LDdCwAqSyB1svZ24vh2v9w2i1/xiuxLSc1pnlWOWUcWdn/KoE/G+TiVPsn
ZmuuXrDw6ID/3YU3hNvoQxbeYq0a37ZGCnRdg/h9PiekhD6q/mAMm4koU7O2ks2wnony8Qz8m8rM
evAQJLNVok4QKDnOg7ys/fwGiG5EkjYRPPg06iOUH8DOkar1EqSISwHHGf2B15HBbawhI3fZw2tf
OtLI8Eb1yajhnOHI06OAoGAQJ935OZaOihxI9uMgXfwYTI/BikUri+VWa7vZFSkxEc90bAWLFkVJ
BdC123XhpElAkRFkNBq1AjV7fiouiQfuOfN/PwtIDyvVKVVJDXUh7xOaIGdIGitVt6a4Mh3J9QY8
FMlRD8ymVTXzOubPUiICC4i26ayNuFTnUhOn2H0+etTkSqvDalBJ9b55w0bbLJdsVBSnCWSH7TjJ
20qYzdtUmgYS4m3fVDBD/QbB9qTELv+iURBlxnhdT+b06IUKOoo2YH8GZdoJJAVqMOTgQipp908c
Rp4k+TUQfVeCG349gmJW25Yq5BZJaVEuFEFrkw2toX1oSq2AMpsP1vwRmCU/Sch/nNpW8nBQS73Z
ca3PDofMlfN3vLoh2wgpRc2m0W68ifqxVPAhWO865ouLElBIj1kVnkWnwYgKVLysP2/NY5h/gSRK
oNbyj9GoE634bdyjX0m/IoiQ4sqWBxLeWwM7zbnDCSxjtJzrH314flUSGvEdQUaKC6pU/GxylzTD
LGXbZ2JooyTrE0eQ32Y5YpgaU9849SEoOwW9+l/L2F4wgh8Vrj7fbjL8bRZ4qECQL+Urky6V/ZNJ
4OA8hxtLZwYydltx0dLvMctwwm7UbJx/Te1AnTttpDsrNXynUFXRMdI0Guu4Li7kBAipkV9Ww416
4qz6gvFrARWxXqVy8rTrp4/a3sVhsI/CAIFztQn3nmZvhCCJ3nD3WekgZ+7DmySNlRzev5KfWdHj
EsPfSNnCLytfbQ36kOFBCMH7Fz0Im2DE67ALzTQypraLLh6cuAsPPSOOiANrzif0UWN1jMzZ5Hvu
6+5yuUVR3goflG5u/CfPZdX5hTgHU2k3BrcrYk46OTQk/2lh+UcHAVpzRgwgVmyebyTF6+T/CPbl
fnXge5aXtFp/69r0w6gO002TBc7tthrUN/t+9BhYWclM7OA4rjNBbmZqxs7m2fYf9dlQA+UtDYs4
XXXOS6bfD/GTS/KZI56XmOfzRzZs3/NjA82RQIBBQSiov0sWVsq09+WNJH+bDT/+aZ6LU2usH2xV
3VUXNdzsFhZqSjDRntQHz/DHudcb6tA5TxFlgn/R8vm3JICI5BqEWYt2xgOoiMWlKkBG5ZkRnFQ6
vKFMxZmesuP0O+spguoZBLl3qfURpJj3tw5je1WRJIadIHm4u8BbWIEtid31PPXssmtBEo2cwEEk
1P1n0YhpHV8zF51VXA2x6tJ4BIK0y0/L/VQhXb8CDJZTH4UZTMcRpciQ1RERXziWXqBdYFbp+bj2
mQ9X8AhqVEYT6sN+dtwVt7I15nHjQAYvl8kJnL2HGnXbbu4txD41xYjByVXSvYJANjaeX57OZAjI
6crW1t+qGIlvzzKugPbdqlMaryiogOd/QjwWpiOkAiSdKpat03P/GzZP735u/XGfiKJeFaCdZ1OB
MxqVdnFUK4xbuXpT01BPDCaQh9yRFA/fDd9EG0aIAzB929YJGzFTEKmBdZI6iLTOnJkMYG7nstMt
+79lVKhgPdmnTVmtshNbU4AqH9yuy9gGOn0MgNfOIx60khF3ZJ+04+Ci0w+Fm68x22YVm7qaqWGU
Enk1PHUCy/YoKE6rtknFEPzLltdQ8419+IpfIWxDg0vCSS9OMmc7kctN96z/5DRuIwZSovWSeN1L
WLlFX7LrHpkjrDh/KGrH5HoYrWGBKpXC0hGF1JVMcJLpbY/ta0S7FX2YJ/re05vWpcodGiC1GWmq
L66VD45CJPYhoJfd1M4CYFNvZNlK1TZLSgYzr4xdgUH3+IUiOZsrIXPcAdUmZG4JYBK+KTdvhwOB
DiI8xbVXgp4oBIj8KeWb1bMv5PJl6c/Bg4QHc2Roi3C3EBdnXMdcBN1yhKnCEYhbBVb+7Um6aCZq
A/VFTPmzVn9/otGdZ6Txcfy3mjHfjNB9wngxD4HYn46hJHEI72e36VXrBTnazE1kBnjF3q/Cbc5C
EO3bR3v0FzFIVD776u1+i9WwHHgBoF6L7LA79wmrkUA0Laty3ICj0GNW9ZqYkDyKJoARvG1DTcvO
TYa8g85lXxGVgplu7uYi8bjNAcicsl/MgnyIos6H/iX8UPMmj/YZ91qYijLfZVV1wfNhZPjqrydq
EcMvg05IQWOEbD8CQjuxox0DPwD7ZXUHW0YRrMfheYwonCnp81EtNYuYnnt+s4fbq3ryyNJVSMbD
m1GMrN495DGKzDzOnfD6wrAt1i8evvRdaIb+CnIcEcTno3WHOGr//Ad+SJjvDkxigYBxqsc8FClq
M+njVPjZ/HFl9K3OetNmnjYNXeps4sHyjUL3FE20uuxGfeRNxq/pRqEOO6ga4i7r2mqNBmQSSxTN
Zi98uJge18H0u1T5lLOPtNF0twDx8NoggepiGeyaIo0YRY+aUdSgiy5qs0sLQLt+Yg+/IAKu4HdC
/mRvRtHUyC24R/ZA6VV/6T6Pl+Z4WBvjAGg4go9w27Aq5VvBBhsWhKwgHVRyysYWafIGc0/Illr8
k0uI8y02/n6hwIWZsAz3zcwwC0eAIWsPWfkqzWajLzBJwvsZ2BVcHCmxT2I5JxL+wA6tQV4mB+mp
/XYXAXrnED7fbqw7bVyZFQkS0SrdTYW56DaQEo8oFDXn5hR6fcNZ8il3EoTZ8UzESDT1Vd0RVDsi
wU72CRmEWfL5jaH1O5BzzdfdZXGGH+EQZSnQA7dQrEqjmXaRRbwzpDcF4V9I/ddZTnzxkG1bKszM
QIzBagtxn0VlVkRV/5J8nJSOvsTEI4Dggv8iKkgvtYGh8Ia35XSCL6vPLCIgAunKWByV1Zc9l6tu
kGm/8B+exGBGjGuwlP860QV0LEj632cJLj5vKVG7Eb1lNFUGGlbPyNU9wFHQ44T/vHC4MH2a4o+u
Up2W1VxFmRtCSd6OY3EBRygcMdMh1LlGgiRdjNN6ZJfFD1Ge3+D1ZD3hIOx72haSdgTlt+uGNBQc
nR7YXg32Y2m/lzmSwox1874Yagae67L9hoKQssdDazhidewymFmQysaY544CdXuTL4pOxprJ6/Bb
JutbjBOCgYUOP6L7WGp98trQJ0CFAX7xs/qb64rmYgVcZNF5hMdGcyH7Ann/3aR/LqOyDXLHQcAW
qtsVJFEr4yZn348EfJBbkRU/KUDkBgY0RT7HJVVnStRxwixiG4BjtR0ASbCDf5p+M6UiUdzpNkvG
+Y+fA5FVZFoSuAqGh1WFqID1OF0nortG5OL9V1Qfu4t7Tit7Vcg6mMR0qG92SbC+faDCM/8u+Zm6
XSDUAX9mpCGiUODUcKkBzCr7g7R2iIPZngZ52U99sgqEV4NjCwp/43NYNIjzyY+KIZ9RbahGLE9x
fV12y+ZkXSlaPX6qG8IwPaiRhbtD/kzuzzXe5T8FPTb9ZoMvidJVOrM4aSbVCx0ivQPAoWqEH51J
0N+UjJqbxB4vr1HZoHVdbLG1I2qeb54Bd2ZEbH5XPoi+zLWt59PwqR0feyitCQlcD/nvJwCIfODT
zlXGtcVTgRytNV+qV0xNwJ/1u0sOFbxH+KsEPYjqVZwh6KLKJhbUsDaf35+RleABhWNqesfMy62x
J+Fj6c7rzrgKktgzMhk/PkqgF5+rqdEI+y45uhvsYqfeRkh+f5wS2wMBAKR1c0Pyh/fDVkoh309c
ot7ATMQEu2S/VfGzQ17w1frjSEoJWpFXd8uH61biBmZGfDLsNsiggwYYSpr+lIebmhI1ub+PmBE7
MpZoQVgNlb4lv3KfC3U1xrldSZVibWU3AXjvzAQ/hKqdsWEGxJ3BCaA5VnuWQciDucEsGJY9AUcM
Vp8gCkDkXSkGs3ay5krP4iw8GZBPbMupHPyzUk564ydnwGJ83hmAqAdzE8cbzj3Vur5y55nxK3Oi
GJoCVFMnMG/z+J2s6WAcuzS6V5owazk/JLdY4BFg66ZYbXfAaSSE/zqpo7+4pWtaxrWK/UnnD2id
wZRgulLlromYZQV8PsBEuvCQDRO83XmTR6RirxGvPJ5CsfT6is9f2XykO6w4fynXbujg7ailckRq
4s1dJhcXVWraVlTQWqc6I55RkR+8xfjgPAwfINdr7zWhZ2DFOjZZnhTXis5uKCn9MjCue3RfIfRo
D9SUNHcmozuN42aTN1wg9a/i+OWIukkHUkta4xK69bsWdKhtqDmm2T7BlGf0HB1ekpGdvQnVsZOq
GAJTNmkUXZts1U8lQ8ZhEHrPtFK4KyfgrVE1arLiXgmzGPaRVq81S5sjiYIy6PJXJKJ4uzCY0Uyt
MV2WguuXfei8lzDTJiUNf7AYQHjBlRWH+stTVvT5WkJ5cKDl1wwo4kLBIqgUbvBrr22OSX8QYVoc
l9qVL9i0AJ8awD4QLjnzjVWVqr7Fo4Djb1e43waIeWrOb+NZ/86ioz10WyfjKjcmE/3JBk0RCCjI
TJwl3b37mmOy4z2IwUmiBx2vKVI+/UPQV3hGTYDPqKhgajREHudIW8kxvPF9hS8E8dCLfbCY9ZGM
pNIR9dsdz/S6zljivmnWodX+Vs6IiF51zTcX5ub1aI/oWtsepSQ86opG/jMdlGgnR9aKWeAp18Hz
vEPHulrbot4RVfnter1+FTDg+I+XS7D7ui+tEn7d873XtlMcPG9vzRncP2Yo8fFJ+RUFUy2dBX4+
jdDJFjT7RtqdysnAUoP/MULArEwFqoGLWa9zLTvlEUNfqECsCoW439OXUZht+/GjfzCriEU7rWYx
on63AHjnIdxgTIs/U0sDEIs9tdp/Ht15E3m9eTBNT0+qbKalwyYFuxpQp0uOq26J6zsnrvMjYxPH
Tu0I4fHU61rzFL9aWSOCXLQXjrjdcUy7JVJbWXWgSPuPE05DYH1+ylEc79Gdmy5ujzdH/4TPrlw8
of3+nxT7FlS5w5IR/m+lfgIq6WYN8BJW+Huow6g52zqCaBXebL4pYmz8EpyoG1SdSSea+2xnD7Ws
FCi3aJQrUbveaLh5zyoOaqmLq921cbo5g5Gn9kIpfrtw38HSddqIeuJFAFHOWW8jloUZ+AdIo2BK
QfKGhaN9DIs1SAD6khj4s1RZzSnBEpaetGEaWNKJ5DbFHfwMfJXK+wiA6Lms5f61rk9UlxXYXl0W
DQ5eq3+u1R9/Cy1tTsmA3HZ3YOvbDkWO9Rh/t+HsjC2OIxrgemdfWgAtfVkkEaZ5h7dNkRvVkuhc
UH7tFv8m/OsH+9b2IDQZuXhTbUUGDKozGFGLZ1VtSMWV3bSXBr6xwFF3rgfXCtjj5P8GKX+IgBRU
99Wen0wG352oAL93kJ0inTWBBXYc2O/ye7JA8op6UMko52SH/J3O+ASGV3dgKQUqkvocROhiUen4
4REQjQULconvdBwCJxuT4uuprWHBA09UAoVrWAv1QM6bTL69tYZKNEPkBxMaiTkSA2HF7SvaeiXe
FIZT5UDxREJGyx1M+guTFT/mkq05s2AZnG78ytUiqACjDppX7GZOP/vPDzrnHahA7fs3hLFl92Uu
pA6AUGXAA6NXi9xvnUfdY/5afXx6GcaWtQhZRhHQIXAOMUuddpLvpwNr3bkJUbUaRkl2/AKtLpRw
q3m7OTOW9uhIh2bbWJEut6RfJjaERLS5jI1q/lUvvT2KeD7cRzyhLNDiMllywg9wZekDPlXUgbQ0
KkByP6cQP7ZZF+52HyzzJuduUw2njP66gQyZ6ANdBkkfaT57DmS61QAWbYqjZU5oRsnf0dCz7yp4
pWTgWvci4bnheTn1r/ihM8yO88ZK0Gll8BRwyxSMAX+C9TbcrPMO79yCl4lLJ3neSbChJu0zAuPW
nBsrQdJNrOZrZIMgWzjJJIGSaQiPGRVGkkdzcPxFZMb7qcUu4qoFbipYfvxFM3CqzMXoAmfmaIWF
6Kj7QeUoYlyEb/kX+onClFW3zN/qNv3SkpT5/nPc6uspq0XOoZ+CJML7tmoypF6TFn51bNGnNIH0
DmHt1U/JVaMt2+8fv+kcPUp7Jnkckhy9lnV+3kCgc6R2/njtkm6SEUt7uJFW7RrHRZl+pHbFab8y
aK6GaMg4Q21NwUYCd+2WBpZ87kfz6suJoLSAetqiad/EB2KGAGOfOlMEyL7Q1ySJ0AfQcMZZPYKp
tIK4q9an4EHs10mCqingFjUfkjdeXixxg147spARBohhDC6ATekaErBCcm+AwUlIC19VGl8QK9nd
DAk3ydt3FkCK8jelxO+QmThyaZkpKPbucNW8S6lPG79GpJCVvaQ2RnnhJMuy7ZPJs2JQQwbmY4zS
d212KsRVLWGf68f4fsgCQ8ywpHFgm9uydANpwdX3Vs1f3ifrInXwUniDIUfAaP5mlgC1b4TMNsGE
ccdMw37sFuxEc4M0HGAiKRLEI2J3OIylIcJ9+KGPyFUQOkALo+zxeUN4yj7xX5K2XcGaqUbcSqmq
h9CtrYCZdEolrY5GFVoo7ZSV+gSGrxvOJdGUCDFRoFp+o2Eno5Ue7XAb2OsXKsGEwU4wWUuJuKlF
3owWORbr7djwIPkSFbfIM95FmRC63ui8rW4D8rkuFl28uoaK1huBT4xrNWjBnxa69mOVQ474Px3e
dc2F0vWzZSUb8n25JFrAl3dDHt6FRVF7KV/ubjlENMlKHUziwCH1+jpP+ZDss6RLxUH9022EVox1
7ZeFYlmRPUR48s7rsB++FmUj2WQJwRWSsF1FyfHYsuyCEtl2O0yXoeXGWh5wdmk5+iu2bkDorbU/
+gAzCkjGpDRhIZW7UQZKINOPyKy2ax2ZN9P9cIQbJrcB2J1gXSuiDYVnhevVPBkTgQAncqOaNYMH
vKwN0Q3U9UPKj6ezm8Kibuz5IEePTNxLrVbP9dTR078mRJ07LJpax/cWL8hFJtBe1pTYSsO1tMN0
qUIvnaMQpzfpV/VVBSSCvqlMX4f1yhyfX6t1ObD8ZTcy/ADd4BECnRMtIGM1RjAe/MALDbvpnlWC
uu0eiSM/RVHOByypqmA9SFRIO0qWlrYjFDVOTMHpFRGdCyr901NoywAKR64L/rt1Fq0CEyFH1eW5
96DS1H3/Bdvzyemygj8Inkw3PHCMo3fwAGRs3+VSPAnE7GE9oTd4Po5/xH2bJpB1mJzVAFnhzzY1
nXtJfb9ZDDLOIJtG043r4iGcdywrPJy3UxnAWNK6LgeAiGTfdBh4xYNq6OPUt5E4DUOgJHZm00ew
Il7R41keV5AWAGdR0xJzO52Pz2BoPz62LzNMr2v5eqj0BkgL1QM/z/HxJ93r8x4C9bJlj51C5yIW
lYnHHJZ9vVyA76Gnc9jh+RD2cdJhPDE+oeT3jpbRJFUB7wmUP9Qs6EoXiG9VKwh7Bc845CA0+qLb
Tr3MP9Oa7ujlo3tkpXWZuNtGHtNw3hPH4zCIYNP1ONBbv2Hyi6SyfgGguP6sA7BfBbxuUJIWAqJV
RVOjtt/koy1VfkJH++0MwdWIMqthAAuvtTOKdpm5h85Vo6H/oPX4qxg8zZSOxhHaVm9ck+SPivPl
MrM9X6TSymCYWZQtq5GOJ9Xogt1Z6tCNGbcNHdxcMOiPG3DbwfjlQgtKQz0ecSsKTCvGigm5Fs9s
RIt9ccaHczuMdrNSqZ/oCqhSeApQdQG99ObgpLHcMZ1NEaK9uCPPoxO3GXciLc9PUCLh4RyNlnNm
E8OLP1865ozS42hipZZ2j8Af81DV1xejcz/MoZqyQJ/XXl89jambCPtoWzIwUeUrydZJ/teZcUcE
wxCwhksx8l1mlf21vjm36G8eGVz3fmKdo9mo3JK0dgHVT4YRzumh7591zAsQHP1OhUHcDkdbKxXV
gUNgdgfqQgpLSXZbho3UtwVgN/ajKORRKgK7sVof2VWmRR2CMGa9as/LNFqTdhlK0XcluTFP2UPS
Z2Gm+mOVVwSfNBm8Gv+a6zuA0v3FH9KX277JfVakaRZWERi0t/JFS4vUNLLbkLe4Gx4HjafbNbu6
h8tbxav0JmUxP8Ixf4vIgWZvD8+ygqiVZCUeUt8zelcIaEZRRsRFZLwxZOBg4LPX9CELIPFJDr+s
BDG/GiOij1Bj5dmSrMtIDg6292TnPi9tAtsEUL4ybkwZ9GESCuiqcMAFb/pYOTKM8k7iUyRi1GvG
0oIlEgJaF5ctNrcHP7+miOTKfKfIa0LB5JMF+AJ6jIWPAaLwHmROOjrZZmvTkAjvqzrb/hbi6Fzy
R9c62pfnKjx+S3ME89OnZhti6XTL8weg0vGd5M7i/OS+K13htgOtGPnc+l6Bb7sQy/X2dFvNv/dT
3dvQsfmuGbATwVIT2YyC3Phvibo2JsgnX8/N3l4MLPEBzq0hY5VwAdV+az5zKcQAW9f3OFoodl5J
k8P1RwS8zbeXnv66LKsDB+4NuG77zRMPgD2FUNMprTLDnk4xjCHzOucxkF05TNxMC6fwYAVJcMh3
8mCaMpjOpeHjfOPcFfZ2oKSGAXmzaZUx0iQ8Ts/qg7unCVzEBtX7wDFPFVtuoz4UcNwIHrT5SdJQ
efCzVDanjRFhiGT8spAzZMGx5d6PzKLGLdOdnfsUWMY/18ghoNAO0uHemWrbU2Z6lFpPdR+do2ON
j2z0dj1SQvtQLlvqv3Aw5ik6AA2FXiJ5hLKel4HDQD7e1G81qLk4jAMqfJz1IQFEvpSHMCgshSMQ
WDYClu7Mz/CmLoqZXsdm/GjrtW7iZqpuftsPTc17iJO2YrdAV9DBJHLz2wGxU6Gt115xnJY2pG6z
JIpR+BOjIF1kUWq/cxZCfYScQMFxyGcymUc5W9DbbohrIFWwRy3Evb0PRYbNpEIbS8MZTxg5Qbbn
O+h7C8VOQtatRIYHCmozuUC0t1qXq4U4g6vcL4retH1rduWYP7OJZV1GaVc/BVkXXo7lnvdg8QqF
X/Dg/Q7faGoUZ2TPFcn4R5PYa80nkF2nKMjt37n4T2fT/K2cf+NMHXZ9xMXcAQTq+sx10LN1MACh
F5cwGAduc1k2n+HYvunvddaOiOUcYZilS9/gCVUYRBx8X04+QdqX10WuexcJ/14IMKEoW4XwsdJa
SSB0vNfk8VEQzTglWB6QGj/UBgajVn4Yl/m4OESG94BwPeg6tHCOEWWKvawk7zxdM6PM0Ao9Jahz
gG0Kt/wm1ihv+09SxAQ10ft2eTWF4zfNjyf4h/NF53/5WcGQxTNuzvverJ6rLmcV0nCpfbVsyDvT
76Xyj8q3s61LDNrl4h8g8b8YQQKDZa1SDu44M3R75x9yJXCcj8pxX1vuGGV0aWO2olHllwIPVVHA
shBcRpTb3UDewb768wO6N9mmq4FTgCLSJwHmqBbwJxZP6Td38jNqY2HOpj8FqJLCnA42nLYoz0SQ
pojVMEBGY1Yc8KQyYR+rR5KXyhamp/2tQMguo8+gPMIZQrvJ7p02FBXNR7oyXe+J6JdZziD0b7A9
8BbRm+rtEkODozH1ZT9zNyNM6cviXISPCH9GJrtTVmZRC/dLWaKowzPpWrQ+uJeb1hCIKiyo65uK
bISime+UPbLWCwpJSzxWvViRyfn2WLh3YYOFdbpVmLufXrLGvhH5duULC3XC0N+4k2htiDMsHOkS
U8NCrU48IJDnS9qF4ish4w5guQMvo31yI8bw58TQsM5Yzeds0xmxY6dR+TGwcdxlOo/aHts51wrF
GunBlGJv8xeCRDwRbnET8OE4ceJ2UySHid13mWADxzR+1v6O30nfcu0BYtzz7/4Sbl9hCuIcAfc/
EI89N+16Tn+QiELL3z73nq0aytEu3CrEMOLGFz4ULgj2ZEGHH8AGTkWkQkmf0gr7a39D1o9OF8E0
ktcuID16UR6CSoGTNA3VOllqwfbDrtLDMCJBQma/gq2A6YbooWLDnsOwO98lkWWNP1L5Tf3YCW7i
/mOsX6I8Ss1OIU/z00HJ0vD8rW9kC5G5NvF5lpA/ZavbB/jeSy0DpVI/vwKVa0kJmSxxgux6Nn9y
wnVkVUwNDYOgM4cfuCNtf/VT8MaN+pt14oTBX0amrDfKKpDv7up1ItfJjAyPcI11UCHm5PDFOTYJ
syPY5V3DU0uwxo58ppE42Ds7PCfyfavcxlLuAqA4Xcpdnxp24xaPtFSH5ZITkWvxwyQp7tlFmrsb
LEIlShBHe3HoGPrNsB2CRmvtur3TE/L75q/zCB1V4cCpwMYndLylTFIvYM3frKFO2m+QHCaGKmUi
MLSqJbP6RXISldVRoLV4sR3s9uTOpgEO0SAm8tVIa6QJQoV8bw466oQeUYkrUtrsAX7j2QeChUvj
CYHtoatO+SgWSUoL3C6CJw6EI5KRl9nKC0wlkIG5kh9oyWqoqao6/TXbM+KQSBNgdguusUUkAaD0
Z4+aVZT6ECsE44vuYtzkg3NwsqWUPoO8p8RYl1AhwFlVL6p6LEeu8emRpdGHsZmi998BEg0sOkfi
HPnlGzyfvsWD7HLm7TPQcqYhZDQs8NdX2Y39Lh824lyuZmCv6rGg1pAIFj7FLVTNa85sVBkKrwj9
f8tyAlNFDrhPaD8K6kkhl2590Jx81WN/9nBLoLSt1wEH5CZMcvqu6OrInfGHZm4N+tSNf2aelS+V
cYp9aEsyAzN7IEXSuJRMvykZRcHVBnc/pAoqhpc7amA9agLFMDW9QjhkWqdvBrqeMqC4IHAwbuTb
9ogJ+ilcywJr7MtseHTc/SBGwsK1Bf3z5WXTJpOyDvuxCkM69iQehFwVragyCs5N+KwlQwbvf8XM
fHnSCK4LHyMomcI24ANsOOWqKmKrVdvIyo7QXzozGVjpptJ9buq3SlzLm6agOVHiQYodfpFRxv8d
sqHcp0yuztpjIF86LjI/AT96u5cs92EYH1DGBZQyMSYR+nmxiUvDVG9Af37hyJ2fVSeI8xPwEZAP
gySjWduOxq7l+1dXjgYRLF6Qlg7z129sgF7bgqriGF9Dbwe/I8tJjKbRuJIlSEa7iEF1fT79hly4
VIuQhx2biA/TEqmeSQuXarTr/g8uVW1BiuYqZpPmETDj3lfzNoTApqeUICqPr+MGjnt6k9qLrSCc
av2uc8EUZ8S+zvjXt+cT/bHdQ2gzHGUGlvoThGMl9MQY25RsAdB7tUl0Ag/nClcoU+QJOLSnWhc3
CsWG3GFgz1TViH6jl/JhWu347YsV7pvDGbBFs46R+2t2hku5oZ9NQLO427RZZLVnqnMLcDjceSJe
OFg+y+TVabxGWZ7+gyYKVLSCZxfWa/LPWrmE61VPet4KWqX0yk0a1LE+UQQBwV5/wRgiO6Wj/A7W
kAGRIgUwEoI4eAPhtMlLZrdWoQ/99Q4inMMPKiHnLXbpB6brmR9/kslsfWf6zHqd8+yhoCaArl6y
La2SS8ajstJHMqGsNBe7iAxuPsL7s6yIJ9EZP7eFeWlw/BEa3PBLlx0K7DGH8z1/piWOPyvdpoGy
r0wcZw1bKItrWtj/NLf7T81ONlmDSbpSHpX1/s486i61GanL04MPqHlDApl0NKnjim7ESpoxfkkJ
UQDg+DZfNuCHL0EiR4QYSZ1zNVLNu/X42DCDMb7FKOSwwg1kHNrjCOqnfOgpge8xj2K021I+KINC
tUocMRjKPixS6V3WDTl2OQV0Ukq7NrAJC9A+ddz5Ii2Tow1NLIhaOxk4+RlOR2sKlDUAfW0lBj53
dupe+Nq42URK1/+/b00qERIVhPMLNFV9reJBDWKAHfF0nWs2ZhdhicPEcNEQ4NDOj7SErNEwGxll
91zYzwZWlRcSOvYYwRgYRUQHsYZi6cA7IPEmGfZdifsAZi1TmJAIHJXsm+7uFsjkqr8DvA7hDk8e
UQp0z1O3RNgxLS9O1s9D0oZX0EKoZmmegwzzZS9YeeNSkuQY58BPf1uiiJDA0jKYUc6voXgf3oDu
qhnGER+VZm/UfxpoIn6RFAVaMFLJMJcuE3959xmL0iZEiPgI8a43c7oAKf4iBbLsNi6c4O/mHFjr
SQElCNMZfzqk31XPgUA2iqT60gHUGVRi6Af0Tx0geegSQNIW37T94oz74CDyUlX8xyEE5xkOagBb
p618Rl5sxW7cxGgt1d/2g8JQKoWaICPfrHgK9aPeqJw/QgRU5qEdH23MfezTUVskAEyFirk3VudF
n/3oeHhHR4Oy+SsmAP/oaYAilzdilxkWXE4Eiq4sVUvIaUXW7uLuWEx9sAaxFLHNA0EpMsYPawdi
ivEO6U1S8ZpmKzLRWQRAjni1SvJVeN4d/krt/16aDsDu22OxhhPNFg9cv1pJUAHNUtwQdN4z6CHh
cxomFxPJVTYKrxxhXEOm4z7ILe0RaSXH5Ly+kOjsSt4z9R28gPz+5sSBO3CzjBeF4MPGcH5O+9Dk
6rpKeWlOxqQAgWQIoKCn3rvD2gTqZcfRlLoF8dXecdTNCk5xcDD1VIBvhy3VK6EQbgNdD7EYGNHL
qh0FkM1z9AyxUU+XUINb0cqCFtRpqwn6aqmwt30fCr9HqbHGqjb+6ZwSQMr/kKPsT6bTqSA7mvT8
5YCeWTM6Jmmccfvq/qhpm7GTRcqdjvisoK9gSNmtxLEY0ajpsuqzrwOkWgL3s9mu8B48D6fKeTUs
QXHCtwkkAZsgsuQVevhZw9gOPzfQK7EGDgnQggQXZB0XfNhhSOsY8BtETvvZKMpEfZuuXTdl3l/1
HWo+XQd+uBqhhiBcCfBM8R0Ky5HyQl1KXijN/L39ooJeEbtjNRNZti+fSmdgnp1JLazH9eheApjk
OlCcrnqzxVZNvNqMf3fD40UtQhDGxLKc2wqMjkRXW6Gevto36j+tQ39gjJR2282ZxwNedVzUJuRI
9MviejeTDkA0yxiQDqhTuxYA0UzvOSu3Rxu7Ppdirp5kETu8jj8V6WSnzVMYrW+TvM6N2OsCwk1r
XX/G+2FyppM0ft+WBfQMra0CY2J9LY/HSqKLOMrXqsO9M60OXdrHQaNIy++gdcA0XTo7yrnMWS7g
pV6DS3AyeEzLUkQLBxrEUe8u7TNpCnFG6jAM3VQ7EIMTob5s/TX376Yk+1OeRb54XOlIrxfIkTF5
rkbLc402mSOH8PZUZzy/kR++GPZh/RA/UGCSwALpq1Eg8gT8WFHseRI3mcpPTlVzMaagH0/NNjVK
F8UDGd+CS8ygYB/Mwz0wKsInJ0KlQnWFBxg/Y+71Ub86MnDhA3uGEPaF2Y5/g+EYYMQBgOiD+4h5
NumPN3SIuLZ29uMl5QtCJh8+wCvzQAcal+LBaPUEoeTfJTMKTj6YkV2fFmQvuq6Ze8AnMOAPzM7f
V25ARRFQSh384f18IqHD5PAvQTwmvO7W/MrNhlt7k7/sJhQjJ1hpFN4p1EVuv4KBlbrDVrFZdd5u
0bFAumRHhwq7AQ7O3xutvOxph9uvF76wXGHg7uvUvnQsCPXw9IDs89dI0W/ZamzQ90GsmAEIFuN1
OQZNsJyN2CdkfPYcJvDGMEu0VSEv8+eCeTKNO4OEUMkMAQsz90rjbr44npbWtY/bK0WxS4EEOL8Z
a9SNf8AHlzjB6KqBBR2zt7uSz799RAMv8yjYSQI8DSUhXQP2w/F43nFWZurIirPA2AIhIEi74E2P
wloqPWCnqDobTwLASlhqRIw426pDh6IZ5zztFujAothRHE9/eWa6rWsImBood9ge2GssnhwXNtbP
wYhddqfaUAeYJHdpG+tLMnaudierfL64N5luFdFqAekhtAiejeQwkKhq00vlYQNo/Ioj+T/7Lq96
pcH+3xEaieqBy5YzLs3B0RKR4djtwBU/WBscC81PE/nphfgqzjAAQr1Xyap9sEVx5rhxIt3F3Cy4
nyzj2tp9gipMd9NfnjgnEySXw8PonOmKHRm3bu1xbnkP893nh6XFJDkd+yBvCSZIdVVuFiXpyiBw
+BxCddJotctZmFne3Bx2SEKrL7HFhNva+4yl86TtVz7NxaoTSMOX/6OJtDF314ORevbQiU4GL9/2
9MRJY7OcT2XhuiYp+yKfZflP9G83ynRBuymmib248Ax+/Cy1sJ7nD9x4S9aiaQtf4ZXFc1xf+Fnk
/pE+hs2lKoChGkFeJwgB/dPZeDXBjpR0pxo4Wtcq8E3f0AneqoNPlvvkYbiHzIuUY52n/vH7N1yS
q2vYs1h59aBh42x3W2Z3ZufZtn/qb3LxqhE3IB/Q7l5y9OlwSS6M0qcjObb5iPWD85+Whwy1qnsc
SJcWz0WSbAyBBc4BNNTWhzNoz8Uykdv04s4AQD+lTGY0SbuKbMbWHcShdb9H5ORxO5/6/l2b+V4H
4Gip/qS5uN08PJxL24YndUqTConu8H+hz8fs1dVZnUVkegadhi0doDBCXEzZ0FgjWT/ilNP8Dic6
OO9LBRIPrySAPEko3kAzO1SonCxDLp2yvm0twz6Bmjh+5ky+WJ+NH2vLlJlvZaUAS1hm100RqTSb
cxYGH2tg7C7FmXC2RLHOyK1YYGgBxZD3tO/TcMyab8P8CDKIOdkB5O5KRxsS4gAQBBbbGWAtNa2F
Emofh6uX9Qeiu1oEQPcJtZaStV3LcRVmy/yCDHwJ+Y5YNOiXb45PoMAwQKI3z+GokEFl/BhpavsC
QjEuWHbc0l4QzE2Hnzrn3c5dM9dPoLXWNQgsXnAx68Nj+5lr7GWLubjJyNoUL0mYHysiqoNDtR9t
evA77P2Xgr+2uDMVQPH+mPnrHwvoW6OFuL8RUqLa+zBqXCM1Vi8gcFJI8iBUtbeJcj2l4tE3cFD3
dL0tomBLwU3Rv0jteTnci5kjw6A8JbhREcZqtHUu8AGF4S3Kl2fVlpU56VdKQbX51Wax/6oY41b6
i8pzrfnoalCjWGkqVGEhukEQAFpLC01zSEaSPNP4TDiNnECcSFh05gRZLi+xIxtykUpXHPYsXJQy
ws3TJWDZUh/fQwlFogmjTetUIPVcNTW56FGvwIjWSnEvF5uJjsgxXdva4lgK0MJ/UTLR7LHE6UpC
55J3eFUFB7/yXIDE01k1qMC0iU8BEzxrAu1EyyAtxXD8TWqcjJvtSQXCJt76uU+87xesWMsZsx73
xLKjxtkYreESqYqHaKOujKxjfD3EC0kaN+NFyv6vcnteqaJ1STBdPWrOz3wt5/6uWygxqJL6WkKJ
eeqkQLfMsfAuNKThjbFCRKjByWbmyiDSCuPTuUcHF4zyCLM3GUwBanGV5Ed/jtlV2RMuQtiSU8yj
ujZ5LJX+UMwtf3Uw/79f3kAzJLPJssUpVl+EktL2rrsM7vAhLz3jZu/HpdIM/z4VuGMXIueFJxgO
ZJncFlxVxvRu+Yhhtj9LR9rM/B+LB0gd4dWncw5Swn7G/mf8uX5C/q2y9meuIHTatl4Odjal9CaL
EdyQWqrubZZHfQ6nvVJOMngR5hjW00xRI0hAA+xmIyTdZpMoi3EeSAct3DKRlXtbWHZdRpr/lDSx
RWka2kJw4xEjwJoyyFcXdWkOAjvkFKlqPDVKIuDMGUi1d9PpKnZKrvN0EGuTkEtdJ/1RFp8BvGaW
Ymf1Rqao1yfGwbDn1n5xB+l/frrIRhzpLQZ6dcXq/Vi70riE9H9XOsqX4860AYZO+7EX6NujcFiM
UwBViweKZ1+TgxbXTUEZmqnUbpNBci+s4Hs8/doaLKaudoJniLH8cfGH2V0FtL9PRS9wLE8kiCTX
EPBNJzHgE9UX/jUwBsZY+s1ChRSKRyyQi5VyRDkUpINjDad5a2hH98Vt5pXWmbfLNKiUV/6wjHRp
xFC1RsZnWQq7svsk6vqvdj6+0QMHcWxvSJDm960+ApoJG9gq49EAZk5T68PSqLHm1VWMxVjZh+WH
gC+etFhqxN+I9fCQCbCOfz2VPb0USOsdTEa1LkEbEJgSRhkNhpQVYiPthOzZWSSNFlNNROlmWOKA
qj9OY7PUeJbhHqFxWlOFGAEVq6iAFsWb5yWwB60PUEgr/bjlO6AGdlk6a4Tv7pwNGlGIvmKA0Map
As4nLBvEDwcU66bsKYEs+Z92RApgxGDMoae1BTBLQaonI6VUvR+eZKlLEaIVfIMehkTtqZQEa17q
KjJl8HjvBjb8+lH61uPZC3UdJpSd+T0ubzs1fCdjU4hvP9xB2yJxy7c4bsGaUcfcACPBlDA24nzk
DbgocPgJHVBWEIpkDmzXpTsYixS8PKECEWORtAHLCKT57bwGqpDuH2yAOdKly0VkylI+amRb73AN
J6YGG5c2lQ5sLWonUaOZnvOLWiKdUpZE2z4NT3McWqvBVqsXMhEnbcKHE/SvVMP+rT57j/Be+KW1
uh+tc+Fp0oYh58w0pQxpHoLoPS38cHas7u6x6YbcKH3dB76Mo+KcmeLjE4Ko9C1GIfzmV4ZxErXz
fCJiTSKj2qzNiTjFNFrin3/G0gXomSLW2iUfmLhNUsZhEomjQOeussLxtRRKYh0rNrfzTjDfTC44
mVcwIj9IqB07461ZA6IYbE+tH45jBWXey6bOmlOnvZz2WTJWHLKGtTiMa8zWiCYDvyM0A7E2WTPQ
gz/qwOEdHuRDE7tNp65Q+2QsdAGEKPvfVpFeTPz0SWtBaxRgO6hKcqyK2bIj4WXVlLxpsCTEz5qG
qbyqQXhjVsl2ABKNB6BxhQ+RSXGFottClW0DsIK60MkycZJtQONB3UsS/VEhIi0U5BX8kIv2sBq+
iK4EIUAaAzNcFKItfzHMlnuHaAuG18w12kmUCo/OvIsMR780udidCVJrjyhTGX4b31xx5IWEwDUF
fGXxwKSALLDkDdS8RHEtbe80zMu+GXsYeRGelmBkOmGd7q8wXh8GbfLQhHEvBfWTqPpUbjh+3bZk
Pa//G9+AEYqmIFYEG7R9UWmIQt4a3mSZ9gJ9U5DMn6R4MgoNa+eoS5gh2psQ2k6GeyqqSSYQQEHZ
q1dusyBrk8h00Sif3ZpodNC4LRsLFHDXcQw9gBN3BaJqEVbH6SkpPtqx2i0R87viJGTD0Qr0WoJ8
kc8zLzrqp5GSAO8yiyxNEwmWKPrn5RhIZcvhSEKjPWkr6Pb3+q2RWCQOIxgyETTA2Kl5FT9HKpCy
7EXPZmopE72p+lQjSmDuwrW8DjioGKQ5VVLA/NT4rFdSFSSFFsX8rkjFFA5f1SNZsk9amoGfBKqp
V3xEQIGH3+CzzYg0diae+3ocrscsZBqAQDRrG3CfvA4VQpYSYEYgQco2mdX+SivEmk8U0p2x0RmJ
vMuDhDICqJWeGbDdLZKIjkZpmY2urWcc6SRM7IwNHL88FplANAFQqc6sfHNpNATDkKEPnoEG+Mtg
sZQhJByBToTCEqg5W+HaS/YV93xDKhwDhXdsIsa/sPrcZ0bj7RkAJZ9oXLB0pAD7+ePAPCzxW2yD
jQK2QvXG8aFHTLYv6PP/iT3MW76QqM0zeAC1M8echSWYsB6PRRqpz8xn0jvBVzUlFX2fCtXZifHS
//Y6JzPuSgV38+/CCZn5A5udYTflNZpCctp2HdH+TNkDIic9F8VOfKKlUgIU4uhcxI+Fa5QuvEmU
th5yLwuBPFzs5H7rbSo6mEDCV7351sKeO+SP8Q8VRcuoeFOsZVgtr402jQStQHqB4rUzli/+dQxK
csnX0txfE2o7t8cOzspVMXkFuG/TOnkRuc3MH292X+I89B04+5YHWyRfbOPXj6Xp6zx71OQgI5uW
uJXXvXyL7xXIpE2a4uIybG7Io10ceAY8ka8tAhfI0RZR0GDlMBDB+7VCLvdfj5bDKDRshReqaQGZ
K4UQcxQyHThGZo661N5jQ13uCHuTHmrsyftnLAezTxdMqL7E4JQ57o09iCDsIJbTpStcSYToI3iE
5E9ZL7mNoZCraEgtG/8fvG2lawegINZqRbocyUkHiylDoVogIBHoY34shuQS3x0WlcEpKRZe7qu1
DclmsfQUiGG3LDHr/8nHEuItkd9Ta7oISe38sLB0dHtPShGzgLYMCFDCQ9MhIr2b5cSMqg/XiCfy
MhZ54ZJBboin2Y4N5kZoVTSYlErpzly9qfAE4WUKDwvMYe3OQMAl0CvFods5lfSnyPPhdpCqIKpH
TZaZ43WvpRj6TMAxl45xNwJwoA7KyfMhcV5k4Eaet/wvjIaQLtc0Xqc/tKTzCP1dmaBPsqb1TZMF
jr3ZKc9nKin8RenbGkdjUbJHRPMkUuqT6NApv3DWMfn4nVhwVUAMl6pPQN8I/vGEzZjdGn0i15fa
zw+4TnTg7Tz7Qt6M9AW6+zbbWHMFe7gOf1I4PpMylbL3sOHsqczSHYrhtrub9hAsaZ2XuuNdA6X4
QJIoazBbPRvPpKe3iFoQoE6LJ9fLGM1QFZCnYLdsKfw99sFXfP4/FYrP31Axpr7mhhU56DZJFn1F
gfj2OM2bqR6zriBd217dtJv8tmBMBkgCVMBErpOCRMJ1ui8YJapzdGtLNsO2v4/+0Da1nXlJZ3A+
D5McYW9YhvyCM2aDS4HXNFnd++ZiM/sZb1NqhnWx7tjecJ1b55baREYcIGG+e+tQqWZsfeYEZxHh
zjLEYHADcc9qt/o427oJqTHqTjBPh/sN3HOIle5fIkfMFnNmWKu7/k0I08Ep/01DY9d0avxIoodt
a/OC2KxU/Zlb4pDL25V7hozOhinucW/M/KeQUiduGLkNUZ3MDIG+amjSAIQ0p7pwuaWE+eKJY4iE
ANPCOJSge1F2EZVqhIGajsQyfguYKpBvFzcWc2XGYn8oDHDRDHo3aJuuSOKQAXSeDhuLVq1pixdD
IJwl6q0oR56AbPUn/aMjdh5VCRSngaAoIbsmHcMxaU4qy2AlLc8MzNFGNV/M3S1MXaeIn03y5A7H
HKDhNxqoYDLGaFEIzDqe+GWSFVjW7ATotvFbydZStO/IORV1IR7GSOG3CrgSrFmoAIPNgszB5Lyu
YAl8KTsHC97wDOV+6ZAY1x7qAXyOQ2tso+Pog0Xgd6MxCegw2bbse35FfX47hsiAoaQg1CLl3RmU
NZeTBSkTqsaimsEJDlX0hBC1EfA2iZM+nWKghNdpluBHA2AL1qsfzIBPilERNNRDB/GO2OWBXTXs
BaXzLP395NuO7oCISL83xUc4rfs5zeFmfnm2JayNM+pNykUDHBfT3qk3tUhd2KlizR/i8duqiQ1B
cffBKjNcYNX5202cWIZx3BCcnxS+uvxynihy9GUe/aDYiR0Tiyp2i+H8tVZVvHiy+yi/9X6P+Cmk
krEP/p8uXIDURzp5jl9S8ZW4eEaLSkC0PS88qt41SqcCfoHa9/RT0rVOKjt8AM8aSTxrb4qdbsip
vCGZrCyGQDrw7lqevZs59jv3PoWsJUSt0/cWqRvo6RHhcSBVvRVvTwKWwuPiADwLcXthupmk+79Z
ACwX9rreBBUPioG0MPjKpR6oN9rQN2SKPlGsVN2PQ3UFVyICHQ/wMwltCvu6wsDYtqrw5a62xRJA
LxFio8UAMw2Bg/xjZ/OaQymYfRJkU2/wcghh/+myjiNb6L98VRNMnWvzh4mlFGReFBnPulIrZBqh
B98bpGJGcCsnyDqZpwHw67fs+8SH9HXJAxkQgDL5tG9pgsI3zl4PfTqIfHi6pO9cUZTMWncipjOa
mTlZsMQeVrCOEeF7/PdB2mbkQGaBTNh4aF+izDUcb3JHGErSL/KcTkdeUrJ+Nv0RowAtwnOWQvjc
n20b86dTC38cJ1xlrV1CR41cIE1j4tZ96TVH+GFOTUv80Yb04aGy1qRVG5wiOdbYId7y9Auustq0
SNAg1Q45tN7KZrpTrbRLzTV8O5m7aUuQxJ/rXtLjHnc3o1EOR16wNFPrrALuTh1pYFVBFYhvNCwI
+JFxpmZnZQZvawOm5s7QRSnU6pONwGfQCjaXPdMaGZFkzqBmjx6g9fi0tcpM63qpRFdjUsT5xI3q
9CYk+78D8unQeRvLRMqNDCFqlJbEUoeNwc28c5b4SJDOBfvj3FBvoh5LqzilSjUIsuGsrPpV53sF
807MC3hoaOjDo7kenPeNvQvET3uUQOLJSfg8ibiE5uLtA/sB3/0aBhzQ9akBIuopm+FOQHiQnq9m
Rdm5JU9mUcxj7AGiA+tAHDT5yxwcTG2jXUEc/C03JL2CsR2MBenKMMWXMeDrkdfogTeD2u0tqqgt
vm7omiUa0BO8u3sOMpepdcjuz14NuWLKC2VkPt+QbiriaXaczzaOuXBE59lxrBFTqWo1PxL2kW2y
r+9VzbyHZHWnuDsLt7Q1NGeNgvIRkAMFGTzB5GSTg7HWBZ2ELjxjIHNZE1RkCmIBeURegU5RRCnR
S3DrnVzA0dOxq+mnAczF62mLAl1wsc0JUHpEXc5PR1B5vmDF+qI16eCjNdDOiqZepvRqmFmhso05
S7qxZovd0DAS/qdrz/l653YrK7osFIim7/ILFn5/VLVSXVuRVcbOYNbc1SqPWTk2LTZY5K8JFotw
5n6Mlj5ug0r9mJjKg0YG3UiE4SY0BtfNDya2p5cy6fB4j0vDDOjyjtJcv7BfMXLqVXLgVCHZyzAj
okWx0wL/JJIL9z/XFil0TvBh0xqvpAoWP4K7QBW2JuaKLAeiJ48eLOINNO5Zx/dckQHXprhTerGV
OwcYIkDFIrfhKWJYLW78a3HS9SG+R4Ukq6rI1OxCR+rHFyzejiGrvU5791A4RY5cSCNrSDqmUYb0
g5neKsvU2Z65JrVxQF2oiJeEycKWHEtyW8gMt0OlDsJhFL37DSbDn9/8UyxoS8TE2wUf/a3TBQgL
VBYQQnq93IrcQw+kR2k1TJGhY5C1DThjGkldNi85it4N/Igt3BYNCRNJ6Ur/g/oOz1VdW9R/vuzB
bOjm3IpK9V4TrlAntV6qO6iAUL3zU+uylhRy1PCbijetnlm4ANaQ8K53C9ib9LEgA+FfaaQ2WahU
2y8PQ6M5OTygE9VlR1qr5Ticv4GtFRvJ4cHTVvZktR6FxrVqVgXls8jhixvX1/y6+gCmkEHjgMrL
CV9dXVj7EQctgIhMKU1aiWaO7jgXI7mho4oI+mnT/SGWsnQpLHrMoDCUmJM54+DO3FVbJqinKy0t
Kt2jj4IHBlL99ploVtNgclV0U+ugA4ym5QcIjJTsgZ29T2/KMFJ+qMvvqSHETH6f2Ec2svPgjcms
qAn7IFX5HdtbqOEoZA02JcY4wErPYCeHSArpSJj48NDndGtgxlW1IZJN1NHOT8PjS7jkNzTnLJOp
4INF9hp1leczw2rU4sKyfI/M6esqnEM1F7lmAJRxJThXaqxJmA/cDFuU9hig7FOkMcpFN2GkuN97
25W4ibG3G3635AD1FgHe8zhZww03BOxUXGsF0tMLXsw2+f7fCchgOVoMxxEpQc9JA1N0vPQgYWVS
xYwY2WCY+2kNCH8SUuLqZXKeL3pkfD+i66/uqgE18mxpKxads10oMdmuA4fn+gTb+gwdfPKBJNYr
XbfppzeTKvA9UmO1uwnBmTcYS3iW79YTlcgunE9k0q9PQ7JHz2W9AtU6bX/5Xnp+bE15BV9rqlRC
xXlRW8wYrD8uhmkaaAL47YeORI4wUkDrTxxjMp93PDm3YE8j8sDlh3DvQ5jyEbdWJPcj0swfgx6w
6Dqy81VVnIhrqGHML7ugx4MlF/Yku9t8x9BOn+tEcEeneqfbCm5L5hAGSAov4VxP3oR4a/xFY+vY
cBnLNWC9EtLICQIxeH8/kpWy0RameaWfyMKvSU2g/1cfSoCqHzkVQ7DscbaBPz+7mS0PlYEK/s/a
twmd+5c4J/l7SYsDhoBfF/F3ijpk+dqzUSFOJjyl4YP+zcl5hcw/XOxul9+nmQmeuVbOcJ03aus2
1GrTNsWA5xSs0MU3HmJ3xX/xJAwb1HNyzD3FcBoKbL/iLMi7NP8b7fzdLHSris8osVuVpN0F/3Iy
DPbryjw5bVZEMfPeulXLr+HlhJ/uj5187b3DNPdJ8+QusC5wmDW3/qZdezwCKCdyf8EpQqkJlgNJ
DqX/ckCnLya3Y+gFklxwBbbNyiCs3+/OyX3Do89HWN4fBIsZWaD2NDJBmDs9kAilqypWzk3uMHC0
AAXgfyTxsE3TRD/5UwHKQCn7IOkEMlgc6+SKqdrEIUdJ6oqBq/fOPOj17D8VA6LgDYGIvPh9ioSF
q9t8SDu2j5aMjmAHgT+Cw8PRK5iF7/WZyqQYO3arBv+F5ig4cAAQEdq5vRpgSH/ETbWvefsoeOj8
2bFNgiM/alx97+68H8/eect3vLl05Q4A0EBpzUDWrxLZ4DXlAhyppxDLUALN3zgyeZ70a69OAyR0
xussqzKI2t9jMdu4ERoy7nAUCIudZzdIj36vU7r02GkgAy0zfUtk9FsZJEgTYj1f3AGB2muYuwjI
uFFXgMOwT03k6u3cUeNxTOw06EqBylFN4k3hkAl0dcoohyU0GiLmznWoeAA+NNQBl6jF3o0KeEi1
8XskNwInyr2FX4/DiIz/2/JXFgQddv9aHMrNh7vcEbUagdaYRJf0QDyZRzo+HabEIBn3eSmnjGi/
hWMb+2wXze+zNy63e/K2vXuJLoa9SLR7uOa6hgOc+9isLEiZTiIY5az/d4CiJo4WvL7iRgO/P0MK
N5pZ9plLJy23334n0v8vfTN/+eFHAXbqhgGlS2QjgomkJTLQKx85fW07jUZRZ12yYB7twAYxY8a6
CJx2XmplPfAIGfBo1pq7eWBOB6XMUb8Zd6jbRgarRx/mWezJvNRfplpmL2Ega9k/HSVLl9lJRPRo
V48bsnUnijBaEjBdsT57J82Z0ealDfDiauo54N/l+Uvh7HB8V2wbHZL5j1Cikl2fx5+daZTsP3p7
6ujuuEJaxh3kLdggppgIwWYRgnAzg3fZBOFBP6vt8k5nxLDwfrVAPUK9rk0tCRhTzAtHliUsQN+U
TokEnpZ3u0QMrg4oCo6B9wqPAJ3xnT3ydu02YkfrAC6GFEjCVtd/4hVDBN8tRpWeovxp4JYvqmRE
RoGFTsF5qFxS6Z8mTqCNoPy8qTFYaGb5cRznKYEimdtP0PmKs06uEBv5Ol73xC8+O5Qdt70Y7TNo
jeZv2X/kZP09ocTYpRevBtphRJgZTJ8v7+SQeuAu6ioLm48BNXNiv4GwObMh3Od7Q5eEdHbUdvaa
vjlWak9uycfYg6LZ98YhrsVvBO2S8801upDfPt+NtPi3n/7FP4SKSp3o0zoDQZh3z7TzEqtUOd8p
I6paB9/hIBuj/lo+6j/iMckQaoyLmS5I/mKD/imTtE9WFxvlgLPJpOyutqJCh385nPTkDRsECC19
WwXR+Fybvcdy6jNX5X3mUI2KB7+J5/RVQg6V3AMzid77Iemg/JfeZS41bzqe05SFLF9eLde/kaM6
lweIXD1sWvgHF2PDlybfFAP4cFRU5g+8qp4P6mO1LrTiJJ3j+IQc40kAcsN39Ma+XDb2IX2BT0Kt
xWmZ78eFrEt/9FkMbJTPIcWQ6338DnnNgoDVfDHjN+7fHnOqgKaYIn4kXhq4KHPm2p36yKvTFyhc
hn/tgQw6nR90f0q2ixr2sTGf+DpF1pI6+i6pSRy7aBu7B6SPFOg0KyYYbxhZT+A0SY8taip6CcXa
UCHTe8rY1gU3xpRLDwYMQ+XwLmQ09jQfBNjTtLcA2vCfuaxobvgqheRLfjA0zymBkA9w1uCpyFBk
pX8KzqKmfVFGIk5iOyatKOIovEPJ8bD8GQEzJjUjjt2DbPBKcORUnfxUjgWKVW9zSYELgZVi/Of0
vnZrwHsve1EJFoMelByu23L3v6NeDcuYymvnPHVYuohVFrcCGg4PvCZ2NpbEhzQCjc4N0UmKtFT+
Me4hjWAc8Ftzbf23GPfO5+hWqxTJtSc5KAQ8ChI/FuJIn1kDvrRwpIlp0Kn/pQVDhtEVsAtXn4hk
vEBPGaryRU/7I5LSTk6/NIVQuVYgvOwxDTQhF+HEc7udw6VWc8X+p+Q9M2ocNAL0sSCQWsTqPv/m
hPECLWTBH2/yawPxZkKpXf5tHyW1FWGlN90EuHcla3FvNVFdNriJPMzc1JZQaUiVj39rwQ1CJf4o
NNmK4xk+gZTUZDJVyKo53nXQZHlhfiL7u5CngxluE12NA5Z/JrZHKGIdhNgkKVw+A8tAeuRsxalU
lWfbrPQjZc4uyPhca7tTckSp+MMJWZOEz9NAJlvvb1NVuVcSj6xDjWJSAJ7ztP/3CPzfmZIkuNKK
+63CnbEUYix7cChUx2loYn6mOmVvmYXPQ4wyfcB04G1ESN12JhUsJZIpEqh2uGFI0elj14UmQGrX
xq+mFhuuEEwSfzHBNnJ6MNuj7hvA80iN9Rfm8Z6/6+FCRtLvzf4L7bNKGgc6pe72Y+8bzmrGHbED
pSRy1qNZ3feB6xT6gDeakZFWfThMKyZTDtldfSQZTlkLKDS/LT/PPQ2uLX/wkNp5tebBjJTz0OjM
VKo++SXSDme8STfeSiL82PuHsxnJ0E8+z27Q1uOKW77N6wk1S1u3xRYzpLhwL7+d+s3KUmBM229A
b/YJ0Ay33A9w0eH9ym6HsHtj+gZ853enxiP1R+9czDtufAJyr1805ftP5XSEyKDC9l6i8964wlzY
MIUG5JDv3nPEV3y8zP3AzVSd/WVaTbBeoGL7dr3JV3KjIhGcxwjvCVAqqNYvC+2/Cm5yt2eXHc6W
h3z+SxWLRs+bm3jvdEut4M1GN47SLiPHzQO0oKfgdgMEkY2CDe4xeMhsZvo7umnLygpAzEBH7C3C
A1oUqifgWB4zhlxLs7XVrVuQ139T4KtL/wFtly0gNO9Yb9lPPt3JU3yGJ8ggIzMHtEryDNuVA4vn
4dgL7HKjcsLEHnTsLaaH0/OzJVN/nK8t09EtVEvCaCMRJUFQd07Ye8XH4Ufoz534NTqRUrcCV1g6
gJkBrTgOuH6t/In5hRhRwfagEv6PUAzI1qzE/tBzAHpengB22QAxv9il/od7yXRt7S7mcypNS0Tl
iL1Ef9wUKdsZ5lUh7I8opPzrp/gOcu9CdHoAN0axuV4c2AlHv/M36rr6R6fWzrMmssTSskQw4X+U
M4WD3tbzfjof5tirIha0R3PKOQde0LG/+ild3pbeu6apb+Pe6ttXT0HLxK3Jft+WDBxpLQCCH9E9
znEWHzyfIW6xy1pRr4pxNgFlTvjEJNw1LWty8nbqXzmXfBIo+NCZP+ObQH1hYG/jn2P04FvIoKZU
78N+9gsy94+jTTeSKdF056gWXkIZHC5paI4+zWwZQXSFlfTw3bRwWRgE+9tuN4Mdutd7X/uUOnvk
JELOi+b3bpU8q0LYxSSvP2fxLx4Y9MVhnb3E7nAFwFGUSMG/4b95s474NeuASFWZo4E01IprYamB
pYQjK2Z5c9XGokpsA9oPCzmBCUHjZXgrAFmh5fhA7+kC2fztGutnQo1qLWKIgNaHpNGeEUrtj8Mw
VSocIhbR4WuUVBVfkS2h37PMSftb3bibqK0Q2Pf4JUSSlGcYDU5mkQAdT8nC2LcI81idR0DoMOJM
2lY3EU7+0haJrjqeWj5sj2JAulzEOMmxZ53xqmLZ08Gk+wix4ZZ1U8jLZPa2z9AN0rqU0LSLwdDt
p3sdJVdu0LvD2i0EHMEFn8qAHw9CpFU1xF0HBYiZlHJJAuLHp8lxvJAidBeCuLmWACMuVXI46sry
5x7gTsniVRMq+55Tk1fu6pUXqxQuI50AtzQC55t6NsE5jv6AH5eW/10xywhBgBVrTMbekpBFaj9a
xCye+C1hfqvsAz1RaEs6PtO0BSkQcAqjUie8zo1kfPz2pc+JKtavwvAusKyDxwrpZ4hjpDiayMjs
AkrE6t+RCWaK7SN6mqeAxtuhcpOn0bjz6FZmczDPLCOk3iushxjUs3t0x7GydprvLmMYGae77QzF
TCSuNKYYUn/RJrbtOH3iO+1phaZ34Elk6xwjioata5ikwUItlTt6qi6Osi4GzIqBYPB9Mmozju1n
tR6t19uBDuy54qeM7oiu7tXPEL/pVtQ//+R51Vt2LtnNsvZh/tylw6zA79dqCOTLodYm5zjW7tWn
/ODnwDhnpW0MlxdCK5AoX3O8ry7frDzAZrWQpaBR38fwiQ3RP38eGsQh833A7OxW8yfQA+7sRySt
UqVaDxH3Oh+to18XbyEg+kyi5BpuGj1T+fByj67QHCE8eEROovf5SOjC8l2B0vAbcVSTNSusHZwX
HnLesbW1c1ZRbRGnGzd8Ltiv1X1zAzuKMj+C052pxNxrg/b1zaG+X6jB30/MfNeRwm5/I+BN40aI
C+mCrD5aK0hjeYzdYiPs0MJJcmEbL5ADG4PGuQ/HV8aAsJcr5G9c0SW5pYZ5/zyVu4auccWQaxXV
UdQvnsd8vCkIl6sBDgqVEXkIdBx/ARRP6BjzxSfKRVw64rcu/JCD/P2gUPj4Cg/hmxtHbyWjWdyr
gzlD/qUaV1qlLOlsib6bcKn7smtK1MCHXHdE3aVMm41wI1HZVQ+qCAzZjgjq675eoNPCh4vufaKl
aCw2Y6WDA1qet1qHGLKEDkE2i7tK3p7pdu7UY+73tb6udEVgbNa+u78ofnnPFti8roIIDNgpS3Fd
yAbm+u0btOUJ2AZNf88BBtyiIQY1gE50YAuXwwLoK/0CvcYCmmHQDpmh7ypX/n0swzxjywcnvEdx
m8arlzEIxnK6qdhchz5ELhuxsidYD+t/D11AJT7pGd4uCqW3wKjc0+WWnz8gVgaxHjEarC0XTXKy
JRvPM1eBaWkXfUTEUIeTlIBqP0/vOlzJkL+jaYuGFvAElf625AOxa9IAx5h8QXrY8PNSiBZ0mN2K
bnPJKesboPDwMuyOWlQNpqDIQ+e7gz8+5A5NX89P0YuUN2RXbBm0HDLPxNQu907G1Vvq8TSsxwzi
Sz1p4St5y12W8x7jgvNgrsXiMOKfL7cFNrBzBkWeJjVH92i9b0A0m4pDWS+A2ozm1h2/l8IDMOLj
KSvIKDsikNmFHsK+aqGtCw3BTs49CZkLfXl0leWvzpMQhfHFmxi6RtrY32sYEOhGu7MX40LpYbAq
pb0QDfQ5+Yl20a9ZUn5EYrXhphWnbdmRzbwCVauBFP64WujUtA/6AIwtiBDzJNjYX3yu18zJRXoC
tMwO0eZBUUIx6n5WfBJzEH7eBlfVhREhslK0IOCyxaqIQ7KD1vr/fJRNVI6vRrR7V96pFyqh5n9f
qEs7u+WbHwj8v2pCRxuZKkS/Fr0FFsMvnOWfnomJ9Cc5l58UiSfl4D9WjC58/6X/DdEjotOR/+mx
TCGcB4z2uQ0EeYC42+Pwlm7a35lUt0kE3+j5jpHbGdInDrBE3/aL0OLYCl7eseSyYYQxlmxrRDY0
Z3/e1DN7RunNbVkr1jKc2H5OoN3pReRn4Vh+ROjHf2IclArnOoLMtVpwdx+f9QssuDNGxX9qjQfh
nm43I1MGY06Qg9yiLpWJGM3SQ1paMx8jvzsaxsb+8g+N9J1CY3A8A+2rgbb08bPzgKWcQjytXInB
F8Qvahf+DzNn3WZoZd6EjkELyWkRKFNvkZ7YNYhVGezn3WJDpnod/Sh7Do3oTr56z8kBfTSn9Rks
gzDssBFc3g1EAf9RtvR66DaN5Nu3KjKYCq5vy78HQOHdJ65/jQ8jBgZSj6r9631IJkyq4yL81Bwz
Sc7xYW12GNgE8qGqC8MIZZGzmQtK826kZUzzx0w/pgZt1IDfy5J262OsiwrWkbrHtSiA+VL8eIO7
q/3ZwKyTexLFkD/gkD36szcfWJNabRJBr1zBlG0qUnymmD6QqZI0dD1LL2io2vPVMDvXxfBF347y
g23xgszzRuhS8RNzXJScfZbR0coMULa0zHoMMKwAvHN9OPQ5teEBTQ2Uwi8Y91udQOpD34eNBJpn
LVKWN3uWEl+/jdz10sdwjXvVb6QpDuZYwFrzf+JDdDpwDbE9f0nHQNFQ3PhVjbbCn3YIJTS4hjOk
ndKd8tUGv6pomt0uiEkyFgFxwuYmtbwrYyV4EQk5SwxEARZUKU9+TAhH1HF1UKJdFs6gAnN5ckGu
bLB25zIgFb/7VLfTXEL5PkciFYMM9kkWgxArBwda3Yi/H6I0J8cmmG3t7OY5tbHrirZ5k8yEwrgW
siK0ibysWuC6ReMb0ripx3CWu//34mF83/jFsSBkryEP+wEGNE7zMc7DPHQJ55CmXWrgMFpX7XuP
jfLjFL5kQMAqkyStxqM+yES4f/g+0glwTyu640YkYXHugcRb0hRSaJ1zVg4iaZUQZtq05BoDNNrv
tuXOsaA50wFaEYXDnDMAGHryxy2qSXZossRym+uyTE97FGf/eF5GHLgdrX0h2tWzvEJEP65fTGwH
AqPGDfpoLNJm3awUA2Z088KcI8KFOqwCNIuUYYgAroAhz1jAFybPI4A7CTkbEAna2SQa/g+q2WyQ
MKZcjCqScspTdNnnGfZmEb9oOwtN2Sc9jVCs1T5H7RIUZHR/8o5ULJmBvO2vu93gtSOMQ7mN6Cgq
PvhJ/l9QxRjwhXkJ7NWuau9sDzk4S6SuqDB+39K6jh/x5oXGB7uaib8KIP4NxQhRq+KUu2swnsIw
9HSUrYSKZu/cigFC260nGuPANd4MLQba1BCh3Zg9k9GK0WGXfbqz4hoZsk2IJe/llxMtfHCmR8Zh
Ox4V+D9OxLAwc6UYqjGQg7DZJQYhKDUEOwoTODP45BpPwRS/Q/EheewfeLpjjlbVimeSzH1Vy73Q
Z2Yf2RiFn9z9ZTjqoJ00rdxHfebjhkB1zzSqnzflI+wEtYd4e0hz9UeUI/6co2XIzBATbXjRnByd
5OJcn1IiWwvqWCF3lNS+qGCkimvHI1VhfYC0JIaSsQuDJIrgoMtPIUy0Wv8dbaqQFj07Z/Xn8rXs
FO/1BoPcMoxTq+1WyaxBRW1+eMUXUY20C3eIZeGzdCqaPvcb92Y1IPE+9SkLbVOUlEXUWPrTbg97
JnA/ltsF0WYTrJ7YZSZ7DskZHE4EpXV2Pm3g3yDp4GVwXY32VOII/gb8Gw8iiUJgvC5dS2TnggBL
W56d0msGitwinyQlOX2bhB+lo8KtIWzOEz5G6w8TUirlgflOPhn7jC/C1eT2s5HJS4ynL24z7qzw
LwBFhaiyKee8kx7HaL6aUaxAoVeCzrpFEZtqhOAZQk2tIlaZ309tcgvhnjmTh9xalyNvX/tG/3XJ
w6s1E41Fjv7i28pG59ICBgaRttywgrHOX4Qg5ao0gFMC32nI3/yPBq15xFgngGxrggG522BvoBY7
NeXgUIiWSpp3QPaPUvnRmmJFULERbIy+aK4tVpxM8fSbW6SQoKqy9WrIhX0qvmYXNVLovR74jfq3
aKLSdvLZymQJyCXd6a5jtEtsynZ/iwkVpatq1hkl7DsOu7nct4qs0guiMrkwDBhBfGBfEMQ7C+P1
Eyn5PrE3GMfle/XldqeEW1bTvvXTct9lxr2mBN+isYK3uNG9mOidAjZs1YJM09gFOKEz5ocoCvOU
2MQxnnEA+c6V8uvwbmSerBHO8uQQ+fMeu057Dplq/V1XbB1aoJVVny/aLfRc4fZaO+XOdnLSkA7c
riANEdwmhyvtsqJssUMotx+R7uMh+mXTfPgM91V0wLdyASbaIIuWauB/velPFYeUhwDilyKKyisn
sUL2gxLqrPCYoSLlf+0Bc1ubKcq5xlmEessSLr8iteR2c3SG/7sahnS7XBWEK3HFG1Jxm5a8P/GO
dCIH5Nts7nF23KIjbgxe6JYbBajni41BFOfYkultERVtfKJORmZ2/Qi5U7kQNV0XppX0nLLADoZt
H04jPT7rXFeX700CYn39n7Kk/mJa98bZBgQ8xEH/46q+a1/5j6Spcc4R/Yn4wp8dB8pkaqVUOuWY
xUC834NysHDxo5IA2zufOSgyvQOwPnNd1pdT9gQaK7BhJfYIGzxOAAKq/GTk3k183Zpj+KS6FtHg
S7kS5PfNOafysIpeM3NWWmN2UqR+Y7Jsw43m3Ans6QVMY7zhK9abyRQzwxGXuWymtOcTo2Q6cbwr
XmjCxcF2rpxAAHe+Yoj1PhP4CkR9VeBmcYxxi6Ky2sapT6NSrRCOw1JZPZhzdzjuroFjhr9y91q+
K21d/iynEmKD+rSaeUUtg6vJbR6BILGaOywLidj3OtMcnG40dW9uu/2zHe/tf5I3ARYe2ejdodY4
o0NtcvY74Fj8r3rxLKbCHHFRhwW2BxNUMvDuMaIxEaKY88l4+Kqo5EXP/IfKFT24MpeQ/lhntV4R
DxT9gBodg/XydjhNuYr0H4aktPcA09XM0d/6oUnrgRXepkJKjpKk3E23kMz6rwVXTsnEgTjYweGv
Y2UsghmVue9xq2p+7XJ8RMPf4PHkIWmLWpy3+wY5pHCIkKmy2bSA2YvzWhYtxkIbFbpCjGAVcQDh
Zo29fiJbXWJU1SLtWi3XQzXzPtg3vksnx4Qp6Jr5DGEsk7n+tICoaav3pXoE+DCAG2z2R53mvLK7
BPUAfZqWgQekb3lQKM/E00FJ1er6l/uZ8e2ugtdlAR2zkNVgQcALmerOKMUUTJ7sROwRwV28M0gT
XrmupYAVRjkz1jOAjH/VaEzlNp9dhhSJWEAuUGNbFGhEtJ6KwUFzd8Ef3YbaKWGzWBJ1HwoK3f0C
7pMHkF5PgXg7tJMC3BlIdcsKzbZLXWEhS/idBiUbdj7s7y3B00Cb9/U4VTExQ3XL3ATl23In5/xt
I4jbuG2fQvfgM/Q0LxKi/Iws1Rg/Xim46GjH0kufVplAJ+xJ6hAx/g1OowiDldzhdzCE3Q8U2sNM
C412k1+Rj3D2byZseFVgJZYn1xzXT2Sf2y65l2Q3SDIXT17FOsRw07+VFCQQXGKnszrvoS+pG/IP
Rv9t0aU092qIOoW5eimBth4xYQT44AqoY3Bx6vMkOQLCfpYNMUQArldJYyLQoDbpbNxZ6+pRjQg/
H9vJ29m5SjE6awEOHCV+XzlIlKf9ixsVUe0pq2lHkiH/ZKfDOhf0MJhINlzU7Dj7cnkasv+f5jPb
cGdT4Rj9KVPWMI6P0C3KZo+63esXT8/rJuMTKkL4Wppa8foJBz5KsN+bcaQD+Q9mgtbH4F/vtRfZ
bGzodf18aEg37PArpjbC6hiepRPBxTBQTKftoVM1SqEYZEPSYukIBQ+tr0jWOgYvsA+rPkaTlcTv
gGVxrNGezMsMeOcicDm1bXgLLT1dBd57CFpgfm3wa5IduVsLH4AC83uLaf4xUVq2aRmx2uPmfXrm
9ftlT0SWED1pVHEs+WBJ+B/RptJ/jtshn8bpMn3+c0SWC1CYLNuA4/7tPp5crqQGVS1yDi5jlneR
i3oey0IlAt9dwf4qxUI3bj9xS7vkZ8f3zCZckrP5Y7v6d6KdJ1JkWsjrWVvwFmRrGxgX0mmhXQa4
kUQuXD2O5biYJ9QSg/69StwtkFkh3co0yQyiEQZ8Q2b/ZJGW2IH3nSYb8n8pYn2AYAStf2xvcdTs
MRdk0UisA7ES5FCAih3aUfsuyQnTTE5Jd3gxDaQ/ZDM2nqeo49gXZglWa05eA3btQqOZPcHyu88y
GVaVarHRzGznC4Ltjj8lCbEGU2ClfAeAJ6wDd4bJ0/553IMndfgeApNW2idZR8N9D6dK13HvwvzW
97NsGMbXgxe0rkI2YlNArsIWNFHwjNoDD5vo/tI5dIP1vQnQiYE78uJA3r1KedntVc9mwsjPxnnH
rSsdb6R6CO+wbxkY20tdue1T6bKGUAb/RuSekkOCA9GEjshWZbRZJ+4kutv98cJuJ9qQOuP2gW5F
Wv8X9OQEMVXeux87LVZTF3Y50gKav7GqRdVWunFmNXY2Kn8Rs9NAq9zpxN52oI6XurboD1/ThPGl
vJVRcbvb5aBv91VgjD9mcth1uwFWLsKfjeXJTxyqVfWT6IRNnt0BGQHXa4bQG2iPvJTQsxHNNEn7
MM12ctSYqi/7HGIKTjgj3nRFd21K6f8dZLcVJd41KZZf7CrV4zYyT4/HfwItU+b1VNUXXYT3wKSs
UMtUrV0SpDzdXsOrypJZFN+Y7Fi3b+WCMBfNt5g/A7Jy5LgRBEmiqGVaq3FFryZej/0HMlLmePIj
BkCdFySdkokWY9ovypeqgw/E8lV9W/Yu5ivZTCBYh0EtWUXYUepkGjOY6driLewjv8iCP0A8sbNa
C2XIGPN824+D5tXIdIayQVWuGSTcWAHDmJyB5jEniyXzkyiOh0a9ZCNjZUwg/wYv2xqLiKaes7Ax
BP6cPEQZOGU2eAkqTSqd0UFetqJeBtmQdoENGV9PKP1fdhkLVd/AZuoPKr53l930RPzUm8wcLuVD
RS+COUctAJCaqd6lCEHvaUEzOLWhaYrW1yZNnteJ9R6tIT1Wu9nzuZs1586bNZAJHTmnjWxYVZx5
W+aWXhxCiS8vRcSPgQplXc7Ql/HUYoBMpqYXhoAKzmIA3d0hLrNWw70WK5XVOigA8NyQh4CYWPgR
vgPde80yNZ95OZI9DsCJDyHs+aJ9yMVy8ChznNQc28Iu3hi4TmzAN3fOJpntM6VPlLs5fMVIzXFJ
CHcu4s+7Ao/w+jvzR/KUID39ltNbqgXN+QLDWwhoY2vHvtx4LRafJOnSQx+i6WSu5tcmlJ61YIOF
DdB+UJgQyw4wFBf0sM2BxGn/eoaQylRD27VqNoRCJhrtvUJAGs3+D17/ZpIHh74Sw88GxFD0SFBz
SVKLOJO7vZSUKwA/d/kLpcg2zSCwEghI5TBfBNGXtdY3o4YXTPfgZwYk//3TqRWgssxraDhQrcBh
F5bIgvXTXR6N1P/1jtBnZvsf9AcErjATYE4o2jKzjACk6UW97yYjBdPOQct6vSUzws4Na0amknOd
CQ6JrFVSwVl5nXVozagFM+o4aHE07EUMeBxKq6Fk1SB2oSy/yKaqvuRgZYdP6NDb+hikcsJ02Zi8
ZfS3Hjy0SCM5CI7/jYnh7NT0u9OJelVjDBLY/sfpFYYezZhHKrWmZdN5FBOAs60NfuP5ce/gkX35
ImE6Qgg0yrnQeVrH3TJ9N+xrWjW1pUoArQYqo4QpYDoaucljCxECmuVdXQXLNEPvuaLymIr+U9zl
yGoFea2KtOOKqRMPYjjVOnHA0pbbFdxQXaLtXTZN5q34IlSEjJbHa0KzSIKlem9TDLdwCwhD+jZK
9UbpaeqeLp5A97o0got4FApgFpPtg9BjxH+2b0ZlYThHpH3lZXFFJ0AMikjYFlaTNLQ3pRfsO2Gn
qTlXWMiu947PsJzHaMzO2Uc58aYvjoZgtteYpg6EccVmEpxmYZz2HeiWi//ACmogFPzGFRVZcNk0
Vpi+15EVplnw1XrxwyR3kMIZlLSm1AyItt9Rg8EvGfDyW5rUJY7Ydl6/VhKHgTXagfn4KyX3Fti1
soZ8w4V4dUx+ufIxFCeWiw78nUHL/6aC9cJ0IYST8eJb5W9faKaubvOLdA5+MMR47thHxrArcBUG
3C5qCzGi/8e0gIcl6DC4QnJAfC0wC+TJ9lAGJ9XWM+c6MID+uC27xjX3baEc8GrZIsCtAJ5otppH
As4+WqOXwoY5yjiwcaZdQv2jXVCbz0NAWTV4qOGxM132xKdZifqWbGkoelMfYl4q+CF8twm0FpQv
+vGAPhwKyMJKc0EgSw2SVSQw+ffZ2/W1I56m1p4w6BaWF7iZ7nRKBtS43fn1HuIwqShZVYuvAIK/
jKI6ud0CeQrvv3XGud7qdVA86qPqboSjgmi7n4YkTeECKFwnQ+i+zXlNN/jWKLpvYZ9EhOKVl9tb
AZEpbCgZmigkAN7QCIOcTfa/4hyHSXg+EVsmtr6Edo2KzIy2ED7Qb/VHRgvT7IQW6mT1t/mr37e8
2U1EGi13Plq6IATEgil5gp53PhlAa6RrFTRCHNN3ndkec9iRyEbBLqqwuhSTQSbNSLowHaW/o+AC
V9HgPWQLfXkvDvh9P6e1RxHtDDJ4EqmtQ8i/MN9waScCwbd7nrUS1kz7jJGlLGn9ncIv5mpK3Vzk
tGUOFur5lyq3MjrcKA+5jIdL3halq8Lm2qufK9IFm4iq7LXsdMek7h/SxZM2oJh0nibwoxpkNiVz
1Hu8a7McOf7+suo7n1LnQUn1kpO9Z+vnHVmFHjshn0K7b3qMvvMNFeWyQ5wFOze6tkoJ9zvFXxOw
47d53FFGtaZJoFgmfFDsSqg5lp3Gu+DnhvlsidiPGXw9mIMIKyUvGFC8oeNObbvz/in1uriZDQPK
0T9Xbcd64fmD+hhCoJ1vv66LhMk5Wrn0ec1z8xZqo6CjImHfli8XVuVezE1WSeDG7SmGSdiOoO+5
Vie7ZXVU66mT5BPE/g0qn1Nm1mIcsKItVVZQ1zWZnJApKoKxrDFxStv+T0/zf+8dRYR2ClL5I4M4
olp7o5V8FjvHev6l7UDyAMnnNNXoRbpbDIOHCnmXvaQ1mjPncEQHweVSXXxJQ9MjCitmz1mkElWg
DIvx51WaZVYemyTyOTLlU/5UG6PixRkRIVGEdufZ6J+z2JXOqa8gWSK/cHD8gEOYcZhAoIMnodGp
Z84t5A/a1nXEXEHe/fy3j5QQKER7fTtDU/uUOBiJ8HFczjbXcghB04mXk4NEuGX3cDlgZda8CF+Z
f/I0g3uGtcBrvn/i23/BGPYTGi2QabbYRD8yLgbLFvMkgPj+Rfadcy/0DVICJwWyFJrtQO2BD+M4
uVKqVjZ47CzILfPBpTlONi91s8YEF21qKH35RFzwlvMMI41c8/9/RYk0MeLXOi2YxtJTPLmPELdH
n0ejJzm5Wcv6KpMvsVsPD2noZLsahe2pKQZo7Hl6/rwG3fMyHmho0hOl5p2E5Y6FfiREWSi3sOPP
cIFI7UsHiL7J6aIY9lDDWCchktLDendQlm7X+3RIax0yyxdMaJ1NSEo2w7E54K/Wgkw4Lfj5znjE
P5D4RbH4AbtXCkirV1R93oVeUDnMf1j9c29JpEx4u5VZEufgDohJ+9Z1NS9skFEo8g/LCbnBozYJ
pBnQC0H11ycg8cSOTIeXLbbmHhoc/XH6QdiHYrdKVp2ZfzNA9swBRQZoSI+yWhz/B0lyt/0eHY4Q
dUMYBM7sbeTN3VKLZwrAQ2ect3musyW7oh5aBzxEOJGBFFhIfJsqedu7XxtLyqP4h6KRWzGoHLzR
l1lixyEW7Omvs9cu5IJJcFdNXTxdYrQLPDA7m7JUOpZeiy2veB9c0XVuBv1ZtWqg3m1xlKr0gL3S
7ltkW9GaZlrKbFMLmPS1u69pjxkBTPtlutncrsmexi1b4S/uTFfxG+Yz5ppWLAwfhUgwOGqIX+7y
cyBY9feeXuBGiIOin5xXfgTNfdlY/jNqpAP5ATCnVK7k7HoK4hF3fZt3jKFEObby8nauIEKSYsm1
zibgucO/6fPW0YgOXGw54jQDkV4Ihz0GSC2Ris1gAk8X/WOYA9KJGhEtWtRBp1PI/wF2yngiWG16
3zh8X68E1fAxhxcJ/D8U83orFHPWvdklPJ3D3uCPPXMJuROYpkx+Q9Lbeb61pEnz26jjHxuJEpdC
tCVVGiLhGWOXqprD8LnmvkOEdFwQimXB+14FRU3rw7vjuuwl21ZLVvnv6yMJBUEBniLpyucGl+KB
ycsLJVQf8st5rnl9dXrDKWsMgGSMcCtcuA2OXAuF23pJz6IqxtFjzmHyPYH3SAvp4V8WDTBscswD
O4vk5gc9Zg6RXm4geSIQl58BH/kWN1JJ+//jQACuTIEfs2c9tEQHox7X0Yajf6UXmKlrjb3pIkPN
0lefKwqx/fhVx3D3CWasOKwWutbPXisjhMgb9V05mEDFrlA2Qa/SvMKxA1mmIImpYsRsiCup8IgT
j/d+7+91VEDoJsSakkls/5mVyBdDA8I9je3OZLJnyU2aSjodzm0+EftnwHWovlsnG/NIRYBkTCv3
WNkRSnOA+QFmaD6vSWeC/qAY/VYxDwNB58psDMY2RTSXcCsoN2B2uAFqBHnuNGZIEgfazLN9aTUU
UfwuTTw2hoCun6i2RA9EHd8fx3vAYY0aRluqxQgnobvNvD3WH6kkvTmWm8tZtfweN0rT04CJBLMs
Pv4kZipjgwlTy5854tRac4pZmLS3hWPOa9kYJef8MBqUXcY2/BVnkxRyLesgpKHBcQo/u8HGmq+7
6s0B+xWo72dvV8/V3SMangKJ84sMTqN6D2NrYd/eW9L+qrssV+YOHQU0/Rl4QaIoe/Iuhj8GxLh1
w5wpNg/rXR4hI/L6egpv3LjfEf4it5tD+keTxdJWlUnpuEtl/Fm2/V22TsacJaSQTEM/I2biqRiV
Z5EPorL+WofVhvycgKrrGbnxeA1ZGxN4pZu/vDK5g+rEkoV9abCiaPd/aARAg01dfRJeQCnpnI3k
fLeU2dl7bfCUFb8w4JM30u1PklTGaykyFOcdO97ACKkRYHZcjZnhdBAM1NrrH/L+/DhtycJc6JVw
jVcII9jzRnEJP5th2alFjeaIUcxAUV/qQZ5ucrQo9RHdBUDqnGl33nEjcS8gGa3ddVLHVfQ19gq5
2G/8aX+x/+6g1cZG03YV4o0a9tgoRIAeHs8kUekQHTmto1KyON+BuG+1BrpFMh/QPVTSzweBGdPN
0Q3THqIMxK6N0IhRbwj/d2GLbgRM+1GNfDWqKA7IWrL4dqxcfNXUntOd6L8XNv6++y5RwZ5DeVOh
NCbYQafmHjonXZ10JFz1z0kQGwW/6tlrwpk3cuCVpNrmPFocS5ui++7VPljqwKcBS9f3mLj9SYkP
/7VltZwT9gU+9CfoDSW9KucT+0jYt5uXNzSXayXco1cpd1tSJz68v+aopSB1in1njekNR4bpYQ3i
eBw0WbAzrpHNM/jWt2lt573xwuPbqc4J7C2lv+96KVw2X4kb2V1q5tZh1U/rWhunlkqTXnT5FRfd
+trUviW4Xi8U37aqpNTM4vThxA4sJa5dMj7+br4EPFivYMNAg3Zh8s2lj/TFE81IIH0vp/gcH5Zp
xtTKZKqUvJwHOQ/UcbcBJqdic0fP+Z+3c//2npExWFzRiM5T5BCbuKTNeBcmy2giEp97osOEVuH1
+ODP94KWHwDuDW2UBY2Y7WxqfHD7xgbVkuFPFser5ct13vwmEcz492nCb9aAr4Gfv32cVaTbA41i
FqwcSCNtGMCRDBjRxz4YKz+OGV8TCDnN2+NQN0MwF739Xn9VWAflfgDqoklbNcezD9GsX4brdgLk
/vwEihta0j3IaCrBNuLliN0ATJqA5K+uyCn2YmPc0i8/0nbOftcZownGzyeNHCe5CR2qlxSMusJN
4GbB6rvGI1keYA+lcoHOmjzZrMV10uHwD8iGvt1+Y9notQmmPV1qwKgWLYxka821NBjBqqtsw4WY
2r/i6rjy+i3xTFTR7zTWqQuqRtbyfCfKz3Y2zz4/GGoAaQSKEf42m35/Qs4hSd9zmgWX3PmwTcSJ
To0jW7mqSwr4QC74ZeBIqITob5RnNQ3N6vMESzMvwJbD1DBcto1n++Lt0Q5FVENP3pVHcRW5+Uav
luQcWQSEE1bKO1qDJqDQD5zmcVArIbI3GZfa/fB/+lkEKDdYaCZhlxLG3Gl2A3tFP5GChrM17Hxa
qa8InkDrUyqnZNJ7OGunE7eQ+oxYbvq5na/VgoNQVi3XqI5shzg3yA/nyVlRfLDAGnZIPJvrXgsF
hv/OUALFNv3I7t8RKJ9a35D+jwl4QkVpWnWPpTB6xXkxoK/qXCKp1bhVsvN5oxJIiVvP2P36U/pG
LEwoFJCtLd+qzgP7ZHA9yls1zkLBmLCx9s3zWVVAd8aaXGfpjtKgxewtfJTr0p4ejWidaI9Ptj4F
zT9uyl44B5bv0uE5XlllFvzKrkXBdTunekAzm43gJcM/I+aoRYhi3/0GwpbFm0Ei4dxUnx58M9ew
fjWaRfmE9XMQmPo6Dko3OmUjkshbzVVwNmrX7G1ACL2r6oYTY7rkYHGxkLMOg8ln/q/uq6zyoIYF
DdaaZeAHuD+YANar2FYM89a5y/xNoCwZWrapquWXOOKhG6tMNdu5CUocDr8E8KVPlNj+0OVHvl4h
V8/3gI7AOEaQZDkyAi1xMTWM2qhk4Bx/G7XT0+GYQhfB5F1RppW0KUzFDRXg8mraXmflyT/Vumyn
7Q2fVrYKkTaNLnMb4vCLizGJyKGtzFlVW75naW5yiHCQNkjIy8vO+Zxw2GNWKrOFoVvSEGHXhTf3
kURD2Xdct7tfOyQRocHbOj2wIpwuIL6xya36MGaEH+sgPYJZLGJ4QDpGFR5mViQlEucxvHWvYzcC
hlm/t7QwEdU0z9UhtYVn2oZNloPc0rE1yGJSNYZiH9izdpX+ML7PY791Yd0tWijVlMAtUXdmBzoz
+NmbTLegDkuKFPKLESgn+Q6qZOsRqV3OJr4ix7/1UILemcXdTSH3FqlFgpxPe3OQhGFMv10Jgiba
pjvekgC3OIrtq+CEaWmVV4qkyyAkJqBgxrp5zZp3R54lu/EZhj6x5cEJWNgbzyUlfxap3LnCbIdR
ncFKygikncjHwjTEGGsvkBu4+HgXzZnipY7CPosXQ9pP5Vc50RlvvyUyhjIx2LmU7c9F1XjDeZty
FedhnbITBjdMGZKJDRYybMFTFFyjAk7jbJHS/nohMgdtrdG9JHvLREM77ZkCl+eT8co9EoPJ1/Rn
9eOaYUnNSiS05Oyf52XcOlj/2VSmRWHR6H1hQmTULLyfdP2l2eFYyzpT9DorTgjS6GxrKA1O5sTt
t1GafOzkLbRLt1K3irzQXhwYuYNBVdXBDj6BUvAUh8KgKrLB/IAXeoMu13N1GMy4Jx+pa7pPGCP5
pGrQBvVc1jCRG95NGtKvrWsPqI69YGhQ2zoG+HIHpXEPF8qK7Je/I15kAdp6tIK5TT9kS0pjRHQx
K6L38gJhKnVqitbcCh9V69vF7F+tR8DdogNZVBml5lYQSIFkb9uyHM/NqhVsINUc0r0148DdszIm
C+8wO+uIXG8d7zlfv9/O+TtzJpSKpTZJCUdOkMs6/+maCunWqasCKGomFUlW1w+9sEm9Ybj5PLtf
SI5xcJRZp4tO/0F0Le9qGJD7GrZVBJJsL9SwciqA2sahTAklitvvum5PgP/RQ0Q/XoGsD4LuS8EC
PDFcQ7yL2KA0AtGMu5wmbvMZnooYqt7/Zuv/d7P6HcxLrVa6EPBwZFIW2SGyG1LvwMEHWqjSazUX
K5ZTTFs80siqvobQRqAHNSp+BzGeGhPlJakMEw4yQULSyVHSwPxqsb5G+a0+iaC0pDtRzIUNR/zy
uuoUcyLa3vEtsGMqQzn8gtdvOnEQLsL1A+oToUXw6l2Txo3EBF0PrcYgBKXxELUJ6ZjfRUrrQdDw
/wFlsNFWMR3c/QQDtbYx0wXBYRm6MTkvEBik3Y43Wh+jc3bnDwRLp3+3uOQoUmIincNjxHaPo1Wc
FXJ842C+xaUFrUC8ArxwGOCd1IT0uDTzI04SwyUtxPsE36wDcPNI46qS9KF/6f4nk6OUgHIGPqAq
f0SvP6gTBxsRdjGm+fBfunCXx/Wxe0YoZEQgABYffOOxmgroqC7hvXHdMb7Ows56F8r4X01anSMK
2n6Z436iQJX5Q2QEJJdMs+o9hO3NCvvtcxjV8neDTsb8zDgQUdNpVfZKwYgtach6qRo/ahF3O050
9i4n6520lrZ+4kNf6xISuuPmvkQn/0XonR2d3+eeVQEGWOoyz8xPdJJKtNNj1XcON1oheD17rYeK
+i6BGf98GgEXxtXlGs5HWmDkVsFckXex/5OlHqRA+7xpqSUSM8GMkr4orYlauwcVlu4HUD5wOUWg
paLbwdi2Lu+laBp0c1PsJFYKLy0JQNK5I1iN9J1kDmnHNt2Y9qg7SakBFicFYFF32v9xNdPCNJFm
njXK3pLOEBC1u7g7SPiovLzh1L3GypWjXeYWf9yZgnk4GtLDPK73L3fwddG0j4gD3Bdorv/efzeK
05ZJfHlCWwHjSDxtyy7BhOP+OU7eZQD8seIo4HrGqtHtsd7C+XK7/jkdnV3nFCZFNzMBICQu07vb
3CXDnebBo7t66USjBaXHRdSOleCDPh4BIGHgc7sGoVOY9RUa19G/VDU41Gnl5XhsgFQaxZRkoyv4
LEWqKkL2ZS1h+zs3GQVo7Gor39l/NnaKvySVLlqfaix3NRGIxStDt8B0L6T6PX58pS8Y0SqFvw0S
ivraBIIlBT/OXNdE9bddIFn2Lkzx9Z8NovxtfjAeu38o6lUwnguJiQp1rCJHw3wvowIcP/xrePrz
Vg75f/r6VUtW8OeLhbxEHjG3vcnGu4fD8wQuaJt0oqeHEcGHRqB1qChJnAS75knbxNhEVBp8v1IE
1IGYzHzAY4fXfre+KBELi5DGv4uUsMRsAZgYLUryR/qNUIWlDUc8j9pCEUwFxjn/bhhoJx0Vusoc
Rb8U4qwoa8fRk0iCoSBLBV9ZK14BTvM7KWWFKjtx0m5YwadcLtUOR5fsm3iQdvscXY2EpogUQAyX
1l0McZ6utRsbOVKrzsWY7Xpt2Kig31VAKcLnIV5eOCua1TidjwYIwqxaHYX8LScHfHJ0MoPF9hC2
b5iaiP9GSRKwwe7gT8teFUzpgL6bHcVndEkonANt340B5brr31gQlWAeNYnXdPes9jnig3ZRKVHK
TmJeXUIB6SlNxn2uG18p3BY4daW6w3xkrABiu00AED2HlWflQkiVojrbHz4y/Wi+9XievPPfAC1g
YQNTA3/+N2Cp9G2Jd65J83h0upVul6AIcqy8Q73/8nNkMaBhpjGwMW3tAGrI2HzUqlOtoXPsrgpN
wz7SBs6TXYKqVQBBY368wlhILrsWmaPnWZyk2U2w9gw3Idgxhbqu6W+91Kfw+p+S3ttWNDaHsAin
Z86vgExPjfVzkLt1r/b89jMa0EA3yC5m/RuBe0tG3H9ka1SmwHSEC5TQnqw6RnyxEFmYX58HxPh7
UUQUG5gwwbSlPJ5ksRRqRwtkbDZ1NRN2/SCfB1DWLhxIl/vHzwbALQ3SYYDl7SJ25d2I5R6zHNMF
qBjKmdoS8oRj6f/T7jxufVqXoIYLdfI7iDT10oMyjP1SnB6NLUu+JiXdBkGAdo3OTlGDrMuTir74
96Bm8D4ohY7FYvbbivgd2vIxld+VkO5xmpFydUqPjOGn1Py2Ls36UbJLMjdANnnO2sVJRBTXvRea
zuo81La5WCgXV1U3Gqah5//gjfUMLV/vBCfLk6lelXw19iSW0E6DzMT4Mue6W+QkstDglsn5RYik
wO4IR86lTgFRsfQKdrg3qk6jCgaOidj6np9RaSbJd29ZFBQ+Im9K1GjH+Nto/liM4cVmpU/DRSoh
o+ZmbFzqhIhecgvdPahc6+1m+v6PUrl2AV91k7TvNoRLy2lL1msDiXUTLDK7UZWxZ8hXy3VrlUke
7m9+1kM5Z/XBP41kF+oGYwp/ycXv7A6Lnrd9nbdCWJqc1+mlp+Ly16MuF6+8oG5D1R/fz8UR52mm
v5x0PBQEz+xL7X0lzGgaLeMpzJlQnswxaf0Ft06/XIOMW4YNVG3+BXSfDmrVYqLAEvigI+LBtk8M
54idZMJkzHohe71iFOm9nSV74tdni93CvPWrbTnL4jHk+LvCkqQhZtzp0lVnzIM3+n4CuLwHKcg6
YJ6O6vhLCUmAS6/r77OxI2a29R5TTVmD9QdwcprA2JmcRR74EvA1so9nSmada2qNHny+RZT5Tdwe
WZ/Ll1GGxcdKkg0eMRiqixqcliPeM2+Wc3Z4agKT94hVlH9hCpRqzlbQeV7alYDn4zdoVlcegK4n
bY7zzqZp1n0Ptskkt5ci6tRv9WZ4e/5rR460Xb9gbn6qKuwGpzTCoZRfZV1nLK8zxbyuqSfDU736
6qg8u1AxcoPFI+0AU4LzgWkT3mqVyvStN7ofn+NArv4XkjVz5r7aeft6imESx5vW2PObYw+t4JHC
VHvgAimentTmFZsF/UZm9Fr4JDoAHF4bRfmNHh7vKbwq8nIdtui+lLwoR+aACFwo94K5OuqFHRAU
+bHs3FN1NFnTzpQh5GWyHLjLxU0uTWDWSbA1A7TXcqeATkE/ptnpqVc7D1bEEHKPqbljno69GA4y
PvXVT8rdtWHNXJ4sfpmUgXuWtvSjVXiimjliRWfjZqEYdwdO5eJP+HFqs3A4sBlAtLPWApNUeNkn
F5D3uEje3oYZzynLebkH4OMCn4WQY47CNnS3nqTmMKgkj+fOoIkTjM6tiKneHW/z7eDbBx/IhyA3
tn+3d1MMhUtfH0T5z8aGg7MtbXOFyIUAE9bEmBJWrYpWaqSSb1PQylyjIMLaOXpLUOYdySQhPBdO
gxYj7fu+3BjbgROfyZxW2asydglAWaUg5deNTi35PXkQT/ZaD/TxezcW8kVly0KxlnyAYb0R4D7h
/6IstKSPq259hErZVjoQA5eZM6XmR9fszdLjter3Q0+7pAK8sPfbITxAaK/SQ+ZdQKapCv61izyW
Iot0IgrKb4TC1IDbGSoBT1TX61rmAR8UFmfQWD1oDuo7FHlJ8CkkqZpafgueZi8cg4+G9zTBuEVw
CZnlh5UVVfbJqBpaTFg35eZvnjNBO/r881n2uJlOUA5Bk8/Sr9/DtbWJo2eCGr30bVvwGSAF71+R
OrfHU/0WE25WOUsehFJxCm1zb4KLZqIqZentyD4tMgz8f4qzuF55iaOPJA3yne9S/s9HHpu7g5hG
IlfwY2zvFGiNu6tpKDJrMzaimNkFKRMaaQhvNovFwhqBaevROuBbgW0AocvFPFFOyok4AMQGvu7p
b7+qfzZJo8HwGzVMJa0yDRREP9jFlQv3UeCO+sin9pvtbT1W/1DZDVI2Cr7UrjfjAeL6AY7vDxnQ
FkvHI5P5FgvGUnULvQVebYqkJMwLfSFgUNZdgb6qonvzOlAY2bPPjzJX//sYz3B4VxsNQbL++Zpq
bX8qYghe2qAti5jsEaXt8CgxLbr1phT3zJbSPopBqRapT5FYwbzGGsIeg9a/nJVf7QJqI56J0sWg
mHRTsLzdAaRpQRfnCSsXflNteoA0W/9zUVs1QzaEAXPIvTR88V5qOIc+WJMP0ZwQGWhZCB5FyycE
Tq0Z1m9c65T+HjdpF2rfki/cyV6uR0d3PdXjLz5TmbByOIbMszTloYMRrhq1grDeY7djUiGthxXu
EaBCOtsmfy6bL1IZZIZbRcN77xXOA0lnwIQYJ7PqaimsUnK/8zWDapRKpybpcRDyfDf23ES+Z3lP
3ZkdXM9PkK8dqOnisnWTcx/mCMHYVqMPuLWrw24601IxfmMGoDgdW8u6fHOiaIRPZdb3UncTAeKY
O+OlEtPpD6c8+TFJW+38gLvKoM9RDxzHByAUsUUlcp4fRAXwgEXBI0mKoq7Hnp9K0s0SMWgqFjxJ
j146M/OoZsdPVsM8YAL4Ot9Y8REuLGG5GRrP3HplkRu4fHxhDJGTzGH2WRrdApX7KrpUNxVLDTFv
V/e/oCHgGtdEVg7MKAq9/R4YElMDbi0AI9QH7wGRU6wspPxQOiie98HBt8Mdx9xhX6W4iI81k4fH
F6q+gCSKe+DQT8mRwOftcpzweByjm37/Z31cabJZyH4ILAY1CH4mSqit80kyhzKFXjvEwTZaYdQh
bqAcEOAV/UeB1Ap5U+wYQoq5EVfm9EXomPKLMa/H146Dl/0aMbMMqcjyeSinU6V0p5K3DKyaR2Jd
Ncsz0vVvqqsVpVJiWBZJJd9H3nIkPEKcMxIydRw0oxDiRSxw5lVXb613rp4idyG3qZUgb4Ca0s5p
XXobCJpS7Z4I4eVC7BBUeVfq0ByVIP7fUZl1ewj5oIhvnGbvAuAqUmsRlB34MQ8Znz9zDo6WWlC8
i1PrkZzTt1eTVse3wy2Bi7jYuhM7acDL04PjaGnh3Yi9KTeRd3Fn/kEdIY0LpJnz7mEQdT0Qat4n
phHEEGDjJA90kGBH2LEL73lqGNpI8Ikw7iqwqteGcQNtbWMOHg/cMa8RCFNwGKGgHGl84u0XvIDz
KwWG0GTg2yB18P0YnVOZnkP9r3RjkiqSIhvsEfvoStyGTbN45EL2+efN1kDLlCUigvIgnYCBGpE+
PLkfC8zx/NRB1e8baWyKE265nFR24bg7QZVwphwLCSA30z5rrntQtSKfJGWOcYCoxnzorU+qeV/J
ubGmWYmRIzu4dTgMOGSv1OyMiWHU68uyXeV/pJd5mbZBJJpACdzYwvkV7YBCsPRCoYzUhpchm2W0
n+ouJ3yLSPjJzCvTjKL3fJuPI6ZQ7eXLD8wSZBf8yPm5FyRpylhd04LBCUkOL31R7CCwNxcEBt17
hEKX8ybe8uTUs38jafJg5AqNVby4vfTMkAzy7y720egikLQTAno1sYZHkCfm6Z5frcvS0+F7i0v7
ifK2vxR7pEa1b3To3nrjryHXxW7hdSLEAd2t6xyK4SYHjzM5t0T7B4v9Mh2KXUIX5cQ5xNHOal1r
MKCkCZcjLoMqIkQg5ypvqzzVzHRVYPSYYUceyRIehqBn0hLlfWnC4dXlFBuH3vJS9hxp3cmHNYD4
quhla76COh1fnYQ9tSGXgcg9qZRD8HUftZeUWtuIisE2UTC18KAIrJtIPxAN6qLv1goL1OKSaqAn
nw32J+6kqS1VnN4SmXtSPJUt6wUpxV/+nn7Ld1sEyrgDgySekHuZ8J+rLMiqVQLZtWdURy5K1ZDL
q6hzO7uMr7Jl+/nZD5X+ZNiQ0E96FqjRyh9HISX7jmflaFqOXbQgYLwzIXY6TsRGwOsYYLcY2XwS
p79ymJ18XtAaqHCqnn1mV2/ZVWHTFYFg0IODwC7gf+St20VnVGt5J64XzGRk3rYesbrCxZEJXdjR
d6HClZnXMLEAkFuNxeJyIAbex4ehFpoktWi5Y5klt6zDOV9aGoEilNmpAgi1JC8mUAGdoVGf8CW2
OmYPn++9P9ihdag6Szh4wMSXI8jQpkI7jWvnkacOS9w5/JEBR1Fg/+abgJLqJOWXNbMghshhcaxN
RDgG4venLTpF1kE33tmv2YH9lF2Akk2pqd0paXOqp269A4gKwE+L+3IDpkTZKPLE3y0nLHCD82eg
xoDbdoMztBaGVjtEnNy2uS06r1K+rgD/fzGcIkAn4y+8g8Yho7BVLjuLDSQj4Q3YJT2dzr1pXmGZ
NNLAmb032cA906/lhV9cv30yS2r7CQfhfbuww5bT2tiplU537r+ew3imWNHR4Am/3TTy/WCuR9hq
k8quCgw+O9dA9YUix8D9Yyra4bkWQRwjLT22o09kVyTPjltmRz7xJPHSrgllw8GVI/Tp95G+aK1h
RPU8EVbyO9TnAVmc4DQfS2lnVmACZsDGfiJxc0TA5dUVYGzO1LaiRTnZy5mPphI4B3nFUCPAdTPF
3okPKMvo5z2hQWF9UFRJVobW9d2Ts6RI/0g1U60LOYGYQu4xnskrBm0pf0q89kTBgu8gWl+9y/o2
cYybE6Ek9uUqNIz3UgxuwQU5hFix9XnwWaG48OpOyP3aTavGlMFCFdGmBZoMGogi28HmVhHfPi9P
QnoWhF0jeXHGvE8C6IDbfRdwb52gpcCTKnEl4vFbk4+YwczIe1U7DtpCGMBLPwcZqmsrDxEpl8fw
flJPyhOcSoZp5MH73a+qTFF+suyR+Q0G9ARsR/+Ug4GJX3bHNey6wwkHu/dCXPCF5c15nnm6RGEI
vX4/MMPpTOrNcLBJq9lPPEaZi2h058QNNYArI/66+edn3AbcSh18Bx/cv9VO0ywnQB2M88ayXvbp
f/+yz8Fc/JWvEgQgkbvWGpRRfeO4P6Wf+1zNZQNn/JYHawe2CUDdyNFkJuAtQ6kwntdOavrur4oX
ReDFzAmkpMv8DV7Br6iOrpXukdJuoD2+DuEg472St0Ee85m2+YuUflkQ77A8sswiZfyx5AE7pxKy
hs1wI+9Em+aHYMLtP3UJ1aaF7Gm4xb98URk9QkvivAeMWS/9JkNhBVugNPFCFVZQHePqEgU5w2RL
7Y0altzZ+PfnSm+4QEpxGdhvpBkxOo7alRWaxbAEOIaiUMy6/eqyq3G7L0qtU2aXWM0/d6lMokoi
WkdmON/nE/ODjcMPjQeIWUZMJs9KGJWvuD5uYXqBIJeSNaKz1jlzU0rMr3wYKbzAygku8Xy0XARg
2mxtD/zFjlTlH+7PILS+CnrdpSmsZbwUSa4tPRLYv+cxz65Y7HxGZdq81OkmbjZNOe2fgSJ9i6DI
gLarKZBFTyEF1xtrvAtqXVaO4Ns/J6jX1r/dMlZX565gQfRmWEsSYtv8HIm0NI+gIJR+BBEdDc+X
rz2U0is1DbOT7KQ4cUMoftSVKiPpsSW0l9iBeiJuGH9hco73EUfIEFQiNdJu+9hLhJJBRzkVCKe4
vKh7wWptCilwW+h11yAXa/dJrRLoNVze4iXGHf+MDggjV+xfEWHfKRRShUYTII4dqart3vWmzFVz
37Ybp1G12BS1GPhwQM5uvvI2Fg6N4ff6KBjGqWV8zmujdW7OU6RsL0s7bOehf37AlqUeGjbs8BQT
02cWa2J3W01bq5LMFkYNfdiiN8KfrtHacvk5Arq+TihErDZUFqIfZMJu45oO7hmmIarSJepKn7f1
s6gdSCanfyLrNGN03nXLPFK5aviNUJUnTuyH+ciBrNMjRjfhF1oFHChuRgRptEgyOwYdS3DJGRmn
v8DcDyCIw5i/cx+6BvE+O8wphLDpifYJM11LgKxcVWbz04wcjFKqE1f8quBtuYXo04UTuKZHVE4p
nfJhXQReqFecN/AOssUcT05MhK3NHK9zMdCTT8EWpkDAGFbVGxkhJ/ahy53D3bfKnSKfV9nFfssQ
VLwPaoyqgo3PODV94fkSL1JFoaLa4s4faoPCGtPn+64A3fQddSxZ2ZHq7sYq+zQlEblBG8b7T4cz
8DXlqadaM/RUObK+TcvKuOiDT0nGhAvdG/30g7TDzB0VVHQWuoDcBfRHui6yFdfuEV5sJQkbjBYk
4ewUO8LVQzs+K+FpZrBbtCmWFvme095BRKc9OXVhc/mW/mPscWoZmMXD4IrB5dpAEI5AbwdoK+XD
Nd8xtH8cf/ESis8wF4G08Yqnuafgce9DUdjtEdpytm7u7NoIJ5OdUegKbrgLCkQZhYcnKllImOyL
arHwDHe60aLUzgrUX5DhpDmkCMHczMEq7kDREkW+jJPGlJe5pL9gQIx0NLg9mzS33Nj96gkBYPfk
Idupf5584CP8pToGBIMQxBWM3aW2p3/aYO23Sa/U0FtSib1LaMfk4I1Vi8ZEPi7SieCWl5omoy5f
LfVLfwjOnU+kq1aH4hFFCvg2r1CHmn7aix1cVhjPJPvIu/cYw34tasFJx+tnrtaJCum3PczNDumI
Npl9J2DHFrXXr/HQM2viEX+KxndDdq7q4KL35Bg4Z0nOZQeK/WNlqyzBgIR4hSVqENKK603qH3oc
cfinTExHq9h9o4CapLXoPDK+ODIAqEVziJ6xw+3Hiur1qBrfJaihbGrZzJ/ezLqXVsLLOAPxX5Rz
bQxHHBwg1fSA9uJyZkP4FBzm2ZQNNF9FET2/wqZQqpUqzuH4PFHmj/zJvN0gCPAVBPsdj/3UaPy+
nFGv3Y7BPkGX6ypa4Dwp1WCMqaPQift2Y+hhy3r5UyTxjee/SnGK6nACqgY+tgzVLpBV9smhuH+A
IEM/YLmBuViGtsm0I6pfb+/uPaL7esd04vAVL+DO3v40Z2YKDTzh2wWTajBorO2U+pANt630dNW/
lIJurmbRUEk2FzpztYLJbWpfeMFXUkPrSFt3NxPVIEqGIRfvNuKzAl9ofophJ6OYBwBQudROg8Kr
rPHxso2U4RE7kBIazhAUB6LqWyohX/qL8dMrKeGyirq7RPzYHnwVvlRFIN4ltQyRr8M4sRPxoxAs
aZVm+Io/Jgixs7galHKnEv+OpYyBNu68FuEkk21G+R3GxjJo8hKZ7xsQSpGb0BEsMseLkltuqsjn
XY1FVMSc7kN9G8oCv4G3CErDs0gaZFufqRITAUkXCUmC/cjQ6675U2mMqsaKD6cpR4tJKZjjKDD9
MwS+7lKCaAbsWH7e5KEvYGdbJOc1IXpkZTi40yimcnnHSfC81wXSznWIHy/mFAF3PPKGs9aBREtg
ALH+mxYD9v9J1QTXSYLKVKDLxJ4Flj5gYGmGgo1pNunNR6BnluOvaDCVfFjZZ0cPiSOQX94pZCRf
t2vxUhGxSn4amdFeThMnOM2V4J5dpGvVS8mzV8zKI1KN49f6shAvQcvNtNDVarHgsFZcUsHKC3xo
0Gn+41bPhbBnMYoN25SZBBqL/r5FUIiwRdJ1KP6HE3vSHcoW+EHld/jYvuXbet7gX54xm/9Jn6Hc
03Fw6JldLWFcWz5uDfWbngL3HhD7Ngztu6MIQEA9ezwndWGCHKAnFyEkqJzIqcaxJ7Ylu86e3GbR
NwGjasHTGy7PogZnV/fDFg7k7eg30gjAGZAAPvXaALJiWQ1V1Pi7XNbXL8/076guK8vA9Zjjfdg2
kG5kB/53AFwCkTARtRkRBsGF8ZUDRYmx5mbXKgxbSiWsMCZrskdkCyn1YP8pJ+smpSi1twMb2UT6
0/1SQggRFOO5fSZ6HyEeqrpzO5cZXp7k3k4yqM9ljilODU3Yhm9KFTuHk/uh6TxO7JS49yZe9sc/
KkAq3ulu+AkHauFJLEGQzo2fZ27wSYGFAA59UCQJymtZvKH9f9H3nSzEypUwARexmPIn4sxnQq4o
WZ04sqB038j1F03Oi8v7YaRj9N47oSOxSo5ngtZnURroO8Tvk0BLQje8gQu6IB75zPL6oOKRC5DT
EAVsq37Bnmi584cHGTAflL2hwmVH5NgxqQ9fRUcK75Z9ogNlBtkEKJEGwCNvEhAdJPza6YsN5I4r
1AVpOqjiYIj3g8cKQ0YZmq99pNUVCNbmGOM8Ue6/VyN0p2RxN79reYNZrVryCeYt0Mwfi9r9HuET
oGhiDG0RcgXHqR9w/vEMQx8PUPnUlRU5x0FIFe0fTvKJs6j4MmpTh9W+YqTlTPSrO6CgzVtcaacJ
2l6lziJB3tYLErQekUk2OemLBKOS537YiSdnkCynJH9LsCS/54YAV4Yimnc+qud0xCpNpJ6upyq0
u3IHFvk5wxfl32BP5e9zwyxvMVlmQPhKI4t8LSPvYPvv5YGuUwJy5tZYyGKXPWL+/tmi9vZlcGDe
9pjUbxJOg2TUZRHG0xFRyBPQvWCY12U9yF+duHvURB8M5srokEbVK+mvhV02HAR7tjNSJ/EGpNaB
72Liok+92+X15K8aG4sJH7XD3OVD8g/olYNGOhavDusL99VKKOzUAahSkh9SoDpNUhS0PZAiEafM
AAYdBYEhvEEsVii9MSf2XtbBOlubUQmzLSuP6LzXnIkm1ls5oz+fP269hJ82SsXwzqoZVRTkf2oX
JltTX7pmwItPSTvwrJan0h6ioIMYeDbm4+9y5MsdNwkHzNoLL6yc2tIhvVjrW4NE5k5M+H35LiQy
GlzQBshmF+Ms0+tG0nN0LCtqy+FmD+tVwZ/iIz2DlzhY2U20+NKQl1mUygK5jaskq/u0KePqc29f
qOy3srBUolBgOOxHcUslVeekBBEElorkbaDuqPTBHMZ8VmoAnYjoZytcK6vc1k6c5kICks7xBFd7
C17O/UgJcjNo0zbot+C8EISNaoHnHc+ziikQs9+BLQf4lRwPWNzMQOVpfAvl0bx6shdi5m/hwKKV
04NSkYwCjjaEcAK0PqUecigFTeZoLbQRFJU38NEJdsUM9rZt7sJG8A3UbmfHjqfLuiAkd/YJyhEb
SaKsbhs6dzTAoivTnIZ7PMSQAeO1QPAbKeL8ocjNYFkpHB1+xZdukk4s6elXeINFoJ1q8PGcrIbi
vNpCNEfZGC0bpkJTCW7Yv4YGAfikvo87kM8w43o/FDZoJN55JvAU3eNn/OEz5WRTn/ofIErkRPvo
P7SOxZm51YAeDc5QCHf1ckqEB11ZJkk5tGRTQdCaylnhoaZ+TFlklKwfE1xNMNF6ocV7fiiDFOZg
LPb43+mEtJzNa8r6S/Px4pJ47QP3hheJTxIqn1RP4rSphZ6Z0IRUTSBsdi5uD65fDnZj1dhL3b91
5tVsAThgAnp1dgTlzpNVq+8zJnwtjsl2cBkj6bgGl6jL+xE8MWD+Qhupko1V+uysKSG34bQb4bEL
lYjsiVus0EWsUkfHIHhX7M4Ck3e3ik9brmsp2MV5XysXDrquilmhaBe3SBfYOESADeBz41kmjscc
hrS/u/kJz6NoUqLyopynfSkCUUmEuFnQ+SOC2TT3TltgB5TF0Rj6mcnzJITfb6UdiEsFJwfi5Dcw
XtjFeEIm3b0c5ODSB/NXwC3LtCDx2Pi5bZ2Zm+sJ7sQebumne0Pyyq1RTSgXcNg3NE+xrrTI/IkL
27IAPRH3GOyeOkfBsP3lHfN3uhB55Ei75skoICubRuTt9FgVtMSHMtDVH1htQ+EL5/1CxbXwqu4K
5okgidi1SrxX+cgMZ432NgqK1umSR7Fo/Ogv5L0db8IzozXnN6oJE10q55AM3kT2SxhR3Vgm/TVQ
4SsMFjRyaS+zTaLwR6MZG5mpCSevjaHXvw88ncuCLGXFJQZrMyNXRxwmWlbRoMwH8P3jens6c4dA
W6A4xggFtKK0tbMpcAFhShfPLJP9VK3i/C3sGcPij9HXY8HjP5HSFDjFUw1mlXxbOt37u6lVN5Bj
QddFBeSktx0Tpeva7mzCJ6qsW8l5OgeFPDlKFKWrasvgg+OwKsyce6RkyND+LiOHEzQVsXd67rgL
mMVM4Q6SISwiRpJZeRmdfPDNeH262GhXkjDH80blAhSAlnfQjdKnRzijpvdaWTlytaurCC5ZkxkM
XT5mhIAg07kNmIZ6OPvHb3TFqTPr7F6xgL1OnDVaWooJyCtTjnkvXw8Hp+bzeQSTE1qgQYEu70xu
SBx/XXV9+vomskd15UBMymTev+ntVa0BM1es9j891LOJut6mSaS7tiY5EzSqerpVTQkYW+1oCabB
Om5SwBAAJOGyx/FuWJUJ6x7UgqQX0o1LgCtxaSUyZAk/KHpGDDc3KnM4Efp4aYojAmEYUv6IQ2sb
Syw/9xv/1A5PWgllLU5iEsGUvWSHiTXsYFxq3EDtu4bWObmrdLixPZ1ZF5QGosorYWfBArQjwLxc
3T9vOdDV6Uym4nL8MtoaCaai95yPUMDPYDJhwOetf0pcKrz79Hlmq/ZFH+pyfFSciyY2p8ni7I/Q
velcsPCZNQMEZvI8qg/ty721aTCAqe+aQzfqLjYYK7QELDJfeEahtx2MnlnlTZK3tS7n6xRIhZF7
J7tKAZT0KFNWlbaRmQpaQq39FkyFjuBXs4S9Aw/GqehZrSBqcYSxSSN7vGwabVStVvaIwpTL/lG8
bAq0/9zCDQ8pdjlxcm/+bzADL0w9K7xY8KmNpVrOd9dICfmOgeu0qHSdI39c4FD4CTGKX+z6lGgw
7cIZgotS7xBiMcUNWpWg4cma9Ov0mvCg++noTrO4MwwCLYIxsa+EBBBIXD5kmVXROqhIdnZSHVjS
UH4H5gV9NVsLVGSCI73OhbSlH6tSrYD77zpqs1814PGZ1JuB7Znp444oo3OttQkMuhBavcMoXy0O
Dhnqed2zf4oYaNSzcymYaWPuPhvCK/MnXSufHPp6mPYO+XAqnHsCX4FokTX/pXkHHqp5sHSZK9Ur
Ei+faLcm+wX3wbWGF0i/kygPHUOQA1Hiu9JzLzVPLMFJI72h2BqME9UzG7scuw7dc2k9aHrEM1rl
s7O90T9gPVtX7VZHw0KoIjErXcPGzWFUAE0ySoB5BvMFNzw0h8n2CAExW8T90rtTlevLjSoxGgQU
thzCvbRaYfeMzmgiYxBR9hwYpGI0G1Ycju8gw0ucc8KUhTJvswxJv82nO+Ldmegmtm5wTjFVio6c
XcIVWCEXEddjIyvJBym42l1oLuJPV6ncHdp/JO9I6Awn//pbh3Hc/d/77QsXAM+e4jTLJhPeHSAW
+nuxFim2jzRnYtoJkeHwS7Avt3y6KEtXLs6uSVJE8gkKLiLQn2dFEGwNeheFYO6VsIZbFo0zK64F
2JT2oCY9Z6o6lVuN7lX7DoCfVLg+ot2h5hk0Bewmd5TEBfzebWXPfi/pgQA2w699z6Nx9LRZFI7e
qYEiOZXg3Y7/XwhYl2z511N7F32TGqMUs2PiFHkB6LOLKg0H9ZxCWiyxqd/hTWOxPaADSfxUFMZp
JJgJJbgSBwwA14nsft0I026DQ6p2W7i231+vYtMOQ1Fy7TFI44SDPiB7lBAEjRuSlXv3AXVInFlV
0t6+M3ZRmksCjCNhtHqYlYdkqXme4L3eRnHQ9G8/Dk7IDsLHwzwE6I0SKO7tFnyT5iR2RqrZBYzm
bZAVPXYvLJnba7i7XmaOjlSLZgAn0VS2g80KXVo9GU8s5WbZukvrmtypBsstjaFhzzHGtauqRsc6
4buJqWbeQ1zCwA5qDALClGAs+PJaMVVCm4nCB51h1jalDaWxQ+4ns+Y9veQVpsw52wM4SMJAxEoN
Psx6xccgiHuouNNGS7MbQpRPTKtWPLpxdY96/nDnkXFUigRlp+bKvuqatPLa8wJeYvYoqhwZfBfx
KnkUpx09Q/RcJkkrU9aN/UAs3ULAVASm7RRFvaJNTgl4rubZwJBkaea1WP0Ruqmt3TNa9NP1GWdo
pIfY9hfogyJvfpTQFslHALrWv68r+58ecHZ+eyP756QOoqK0g5yTE8jWaCfxRLY0dpKo82Dhe8Ei
yBfqVoseSwWYo9YK+rWpcdboLIb/K94yTAXgKhmA39pJyXDSTaLhWM56SAmSuEAbf+gB/GiIgEKw
W9P+2YCmUbm4PKOGg2ss1tfGViE7N0eARSUA0awKtKWAoDJW/A3NHwXO5KROluDPVomlHf38Q1Jo
72oS8LFqJ7ehsp6dIp0Fyv6vT4aj7FmeBFeG8puAxb7onj5J5bVCTCCP4c/CWkHzhTJbDwATjKsB
nwfL6e93U634Ov+w/abSvexBRUG89Vw0BdjCbWQVAgG0AWkPNf8pRsPxuBvk5Z5CUn8KyBHggAPz
aDXXfbqs+U2QjVWmpOzpCpk3lO5EAPBPDfTiWnZDvoKZxZvuG9x1ZZHj/CDsrlgALaJfRanPq0Jp
sBDfBXfipq0NIR2crJOlSY9zRN+XnkiF7CAVVx9Rry0l+zY5np5XWfMxa7H0kRCv/CeciTcz9bFc
zO5twCKDAAMMEYtoOq7/On+6xp5WLyoFQ15gdDZTLKVfbOSZZ+3MtCrFnX5S8BDzDmmVDTsT+CE7
ebeJGCCeRhasDMIQf1KI8IIW4GnQDTkJh81MaX0AgCslhf7+aArvy/T7f9FW7ur8Kbsk8Gu1FkCF
nfg4TpQgkzwh5AkVeSLePhRc1CjFcoJEXud5bgfazH7YSoEtv0sUNodjmGoQ9Z4ES1bEzOX7MRs5
A2h2ZNhxecgAskzjDTxBq/AqUI501KaXe4KehsptMRxIXZGgw6nelc2tQL81PTBgX2CGSKSJYGV2
YLf3oBRttApcIE46kzx3YeA4B6L+7maHd9Nxo5ZWNspylfNT1YbbwgkdJhOB1K/KjR4eginCoFV5
OeRjxRwk2VHiW6rKk3vGUMRRrXvVZJ2sT3xTBSS//P+uVj7Jawr3TdJQeF11DXRKK7+5WdpHP4Iy
UN1mTSZMsfgzSLejwU6p+PM/abzG/8HqXo8KT2qyKRlZ8cZAg5ouoKa6xMft/j+C8G/1FrM5VDx+
NHOgEf+5Z1kV4l8hQWBa1QBnCDxYgwcV8CVRpAfvNOdm1hi0Q4qtYm96DUeDoF/yr/T4Ko4/rLxb
R05f2xcQwsKJBXigeh3CnvuNaMsnCLLingApeZmh77xmjgEQPtIV5S7bMMSSpOHhdKd4TftWRVeO
zHQEbk18XFoo+iW9iAVkHPCdlomZvs24LAQryQVNjlNY9RRMBqRi9YYtkD9euu5W7IZNYeU6u53n
Wu4XyLcraI/7Sm3Q8WgKrLZxSr2xPU+gZmvWe2Ltvcha8qcB+1rGI0COPSrY64NARfZzkl5xDouc
08QwoupMOcveIc6h703rJ76nKtrzVyamIep5aA6e1OO8XbMcOnlp13VssONllFEvCKszAO8HJsSW
viYgfJxx4pUan7CrCZiOwV9c5urPYuLES9Wrl1XKa7ap9yNe9zOm2QB8vi1Xrj2hXJGSjoFURNZo
3EUk6v7nKcw+QmgzvEqGhjfGdzJg3YtzTON1FY6/PQmFC1MFwJOh9fu3uadN//YoIXIdg9ZeEcTA
EMn0DwFVGY6eHrcuzMGHCH65gdCI0nP7D/pCLDuslsJRhqbk94oc57+qf1bfG/Bhe1H0NrgwcGoH
EWxgrUSGPch4fYsHr0l/VwspcTt+0TDYgS6axv/eqriFZ7ZWsqyWnRBhhJ3dk8rIBVAtOA8X86LI
Fvf2K0EFU6km7szUEbOuHZBgLoW784bN8SkvJBKHpPXTiYxle4gAW0bI8KVjYmQ7sXiyCc5NI7m7
ZTCCSrqg7sGYFas4Kf9ybrwPA/ZAOdfyboFqRzDEM8OCt1NIV1qcil76lvx3YyoByuTcGy+ABh/5
a4E/FKyB750cQPsoe4NM+MHDn9UNC0dSKVhzNWVmzxLs2lOlHRTJjNZwGLYNpj3g/4RAfB8vay4A
CfPsO+/3wgEeEspQG3vhr/2ygUSHInSw5h9IAA99JQ6B8ORiQT1zj+Mh+seuCETJJz2HOmaV/dS9
PZKUfvsX3omYGjinqNSpYIXMPkRK1HQbDHUjoa2STVXcTs8HOzXpDJS2lKLwDu7ZJoRYtPFM3Gff
rAanO3++GlHU8//v3z3LlxQfwXBNii1jMF+AeVIMiLJwepri6onpe1VeXC08JOeqBfyEwEvpUVPo
UmnmP+z2TYOgjjsAAoPN+yCC1X1WuzYsxfW6LrIyU0Lbz5gb+ZKfW6xGczxaPWzJtIIurPyWZgGq
keOe5BtsdUnyfifLLpoGFR2DSe+0i5RP64IC38HMgzVwSyV1hxHr0r9+gPI/8Sdu/7DZlsOuxfPU
OTuLabXN/5ryCFSa8xcgA/AOb1uMgu0MpD8aHBB/E0WZQHE+oUttBgL0Ss6Qk8xMXJUk3coL/yK5
E7niFm8QP40mWr9N95TiXBGj1d0DFe+MSKgiaesh+3g9jclZQlCgx02TnFYwQVXuRWy1V6NivnVM
H0+ATNynutkUifOei3j6ciVBTjQeM1hoJTevDbPwMQqWXEbgMXqBGYbZucr3q4ZeVnXBcaQMS1cH
GIVC5x/t7OKKIeeEPpYwjJhhL153ykyf3o6BWGEq5ZE2rP+rarPltXjosb/hUmTuWU+/OZEgaUQp
Y9yD8zahebKeS4w6YJpPwGsbUK/1pK6UVf/4GNwi9DnHh0KBF9bo2VFLycWaA8wOmipuZacBv6zs
nbbBVHb74hNh9UOWVc/J7ylnvD9zac7GMVmKI6SxZs5MH2OIry7Yg5TfJ1Dy+enQFFxXYnM5vZjb
PgqQ5Tc8UaHGz2dtL32QuCmeeP3PTp3G0OzElRcJ8b2/VYFoqEBVGnExhfj+Er9RMTilifmt0+0L
+epJNFkpaDXxv5ffDnj1/7HtrnMRStcGzu8x/VRmN2VjtD0y07uyxbbpno8Ck75X+hAyRAWP+/cG
yXY1FRQ1dZtqSOyD6F5I6M7XjDpKTCW4IymkKmGbXBFLNGhdz8NQrLF2q8Ru1eq1VWczWqGqrT90
I6ADFdUHuxUcI3YVkkDnXuq207i8T/M6Hr5lXnT0BEt0ypzLsXu9LWhAnVTNgI2ZHlWMW4MzGvcO
gmSGz697eZZKdJxpV0/Fm9asjkLwywMxO0gMmKExtm+w32eGXX61EhbVbajG2tXynyWcGU6IzWeT
3ua+qN78y9f0Pd2lE2pwyDe8x5Pw47LjNw/z92aHmt3VrdbmXr3krJgz8rEJtYIz/SfTbwVD4po/
U6IbVA+P7z5mBvR3efm2FzOBV4BS4kglVGgiIRLV/v4jD9V+pHig5RfIogDISHFLxqLesbjgC3Mj
8rva1N4wdnuWpVc4/mhMx4tdOu1TDoRZSRBrYhFII814MOPlYkR/bKb/L+h1RMeyc7SjO0g5sPvT
VNRaSkbh3mOphARAU7wnICUXEoSUfTZerXcAFP+EEhcnkpAtlqm8ViSx0O0D9tLtYGUwJT8NVShV
I0IuJ9D8a9tfJiD6FsujuEy7iy7WWwpFghC/1xny/5Tm7Q17bQToOdf+QoDDvU0Mfe2oF3ddTZHG
BUYkj3Y0pszxDEzAKQDrUZShJHxHyhyJpbPb2fZoPOZaVvofJ4KDDpk+IM6o0egIlYG7jRQvwBHe
niSHVZhVJfTe596csQPi3yQxrlZf/bFiw0XDazWhvM7yQjlcJNXZ3J3XGQium60X0xv7atKcUVS/
DmnamI/6qrpWMKwKOmqSbuRQO0VpQsK997a7NyLOzv423mexlv89i0BYAOw9tmfm8Yf/aM0njG23
/txpQqXPScubVf7WmNgo75S8B7F2Ew+HtZ0+tNoTX4kCU0ft35yHZcuZc++/VB2nkzp3qkHbMTyD
zVOTTsuWeAoDeRacEfURBmWjphWMAAQUkXJ88TrxJUNpkojzF1V7cKF2xAxXg6vJTmbQ6pl90sKx
DKnu+sXxmIXdLhQ9GDFq3+9aeknYNF6u0d2OToZvsEf16PB/mf1vm0+p3R5p7nMei7Loyk/4iLR3
QI/SvfRKzgkIf4Bx3iF9W+S5/phfRxdr4P4yyft/MpVqFfu/kkEIwHNxhMhjVdz/+QYNdZrSp3cB
m3FNt/5Oj9P6LLXrcIsKETlY897vy5G+5Ruf08MM3Ku6wwduRCSPTZFK+/qeXI2FQMQfNb+F2+ao
AcuXgEpPi/A6ETjNqRM+dyKj85bDaB3eE3UqCQYEVnObMvmqvk+gNS7sNO1lAXFSKj/K8dDJ3DsF
4wdIUWEV6tNlrmL+10qR7Qy4XAQ0czaBeewFwjcFHEwM1h9dY4qdN34mkEtS3xJbT8P85wf8+k10
F5KqxDIaUrFz7kdj4lOz8w5kjAfUndhIZ+YnMcRzD+b0p67sV5ZF4sJI52emI+etA/r2GXeiPSeW
vtrNrngm1KCP/mG0zfHTtTYZUDp94iFrvmtpLt2+d2qrQExJv6jIiJ0TDi8tLgZH48VAcoT83Spm
LiYLbOyjgHm4YQa2+f08N+6o7aLucwkkFooizXP3LTpx95x8xh75+CLol9Ep6fdKWykST733Gnlz
mZ7qu9qJk7IX+/6CGU06T7eFnYyHR5tYINJrRRCY4AbP5VmI01epuqWi39te3THQCY0J0JU1jCs4
NZuP1KpOdJj9vRFJMqm1ht9XjugBfTr/lgMaRgpd6Hyr+WoOvbf1kXuszFa+p2kyA8wSDmxUqIJc
hYjeqCE3FOPJlgeRC7YmLK/v9CeRSkeM4YFIf6D7MZYGYDK2G+Kfze4RpEHk6mDu/+6MYjNFwf5Z
+tsrdTX0dcx7IihBub5QXhwPBvkzzcx11wLWWZPlab8cn1Tkr4kQX13nXNZSWswY9hsFYpUWM1sD
RU9vkfOyabVWUg7xry3SMPW6dBIQUKMQ5doshYu3ajNggJAyfJrUhxcIMHSlvhYTRn+2iRmYYNKS
vbdsAeymOHhrJN1ljJx0PeHdaSd6DYH4LZ+nfQp/RXhs+YTAxcHTxWZuTdKoMGYTuemZSrrIXQCv
Xrp/+jRdKpDaLGVr8sAnH7jZ2jRbPqPOyfFHrCGeYWwFbEJe+L1ZetXEX4PVO7A54nyJiXhBVtsh
tqxH1o3HCUCrNri4nuswXPJ+gbf5P5tjVpBJRUP1vQ/9ea2YCHWysC/l7IOM4wf4D6kXCk+oL+t8
WIYPLH45az5qsYGVchWgBBfKCQEXBCrWxEng4Vr4GKWUp5g/192mjTiWPgRSwcSpEzm82ADXqDru
hRAT8usjvJ1aryHx5DifMZeqvVaQnfFgIQfPWu/4AdQyCVOiAz0D1tiGAfKFdFgMy8D4uiJSXOxG
wcJIbIgfMFPivk15Y3YYVwx0otbZVlZvkG74gHSvAwx0jhjMLf92ncf8m4wAcoT9SOgrTjH+wZfh
PPBfaowLf9GCSwsGlAyO+I0C7mWVy5spqMN53g6PezdXsQUjxD7jZDVHTGBXO6W5iq++pMrPHeX1
Nzrg+GJNVGBIBacvBcFtQCac7Ob504pDX9m1JHDyHs8PizhDEUql/2gzAFdOvic4aR/wm+Tjjmit
0aKC3O9T0Wa5n2crecD+rtSLq9DX72igIPM3T6LcqQMuC2Tnf/4vcLJdwuVZuETSXwucZ+HmYoIr
JPPFeA+WgTF3QAukuqpq4Cyd+26Ptd8t2p5lP83kv2n3wuBq/pDR/FEa56Ca4XMKhJuHVWM73KeK
w+7azYLQt3m1Bkdc2TJr6wlaK1Nnt8/2tn70m4GRWmYrT5/QN3m01hYlBt0S4K23yIuNto9SAADJ
GT6KPUG+K4YRqYLEx00etGTofVrs3+FO7rDB0N1tIZ5HpDJ/0SUy9yuPRs5He/3ORiL4AB/rom3E
magLulIRBwXpEcB+SXhkDwqC0x+afn8kvTWdWgQz43dmwZWfdXhI4pO+eph5gnsVnP4HtpprkpzX
jcXUtUMfMJI3Rb5Q8VzJok4D5FqzUg3zE6N2hVbmRoD9y1nr+HWSwzY63DEOtRJgY30nJOFXiLMD
JBfOorkxzWLpmNmmOW7iK1DNEcZTsqVUv4evZYIUX/ze+lNr7mLo9P5xTGfmoK7m8IVKY1VVwV+m
KYEs8r5kyc6aWGVsrltOcOm1lQ8FcEz8T+Vgq9jFfhxHYekW2bhLOuf31Lf8Kdfo0MWzT/JlgAAP
zJO8Yv8LLq/e53XTh+AfOQidvR2aMqHsOQpIvkUcGqgfx3iP5nnrWWQ90vg86vV2eDGpp5F8kBQR
WHYpCitAaJO/BRI+omCH07j1wHcMTbaht0GA0vtkadg2lRUE8o9l0kBeYXitWm7mQ44ZJUNGultC
uQ32+cqKW1i/C1wcs4ahSSDvk3DpmOxRI9zAnnL2v1ywHQyY6PbnLkPBijHbSKk1nMvYhgdKT/56
zowEB4Yknne5teYlQ7jDaWwp1H8obkWYKs0U4luHeQuDYpOkKEUBUMdUfORGR8ZY2vo5sBwEvIr/
0bqCS76BZlbb5udXoILwNtCyKSdfp8NY7P9VuIu96x1JfS/KlA8j6XaL/zrrlljeQ0GqEWbkx8q6
fp6219dnUHDiz1AbGFoW/FjHYF5hEnzS0Do1LYnMTpco5jd0JU1613KNIqfDCziTpYrIm+zr3VTd
RUcHlRXi+uc5k6AYgNnEeIry/y/rmSooWliF5vxcr/iS1a/pnj/s9sWoxIMs8pk9SlYx3LWow7c4
irFqt7IBQt26nK2OwyiijUesCa+TJn5J21hIxAY/EhY+5MTcXiZwAz9qa4vLCiUACKo5gk5CFTcr
w7YtD3iGMCi32TtCkkCyiFHm0Lf55L8lGK9SFAxrVRnXuU8eFcCOMwMmHp9m/D7f44FS6QeEhYrw
0TcSojYFJAIBke7MX3Ii/samkqUAjvCFJm2f9iu7GUQR7iOBxt0bD8IBtdYWht7+zIB2yXJtf8Q8
yDYl/98WjvNNlynGyJJfnbqIEO+Sk2Nwwn/lxMCD1bDE5j+yZ7l0sqezr2cUW030+239HXaG7LHx
hsoSZ3NWVXKZxnKnuiNVpVacFJiyC9/1FGRbdsLOLTBFyCzum5BZzziVfcSJf89KOR20WucZupjN
bXCjvAEWXZozi7AI4LWwaLJBDl5cRykCXoYeKRFk7euPRIZS0tdcKeYir0TAXcU8nyOKxN+KX788
DF/zQN2+60TSJTtGE7Crt/vPPNndSkrAW34xxqeoQyJtxFL49gq8N6LNQFPTzaSZwYpFS6Qy2HK2
PGybiZAA82ShCcK+iM86McyAEiSVMHhV7Z0Ty0vYtHd/zoglSt38a1kvnfUlSWLuIye7uRKCVROA
YcWeZnz0tK86Y0Jp8iOLU87D4tOCZrKJFrPCibhlIeR4h19eMlq/+a+6Oh5IpvLeF1KCXHCPjXVD
Id6qyv33BmccWhs+VJQ2tFcnMmcRYqNmRIKKxfVoibRFybpOXrOKqMxRciqMGJQKwSs2Z08ff3TP
LS6Un187BkGRP8KLDqj9A880Sf8eOUVSk49e/ZoxvLFXTpsHESsCS4qHtcCfxPdcdedQ+OQE2DTZ
yHZh7x2oNUVBc+s41hV3k//k0PugzGbJcxbAM71dOtrqnqilspP6Mxch5hHlVAmmKVn1NziWWn24
ZQFmhnplUKuGjKGDgVNfNKDYKp/w6uOFtE7K0k0aARnMaARuO5W8W/YCJrVl43IGghQqW8Hg6NFw
JG3hjdYDGbivEpIW5K4nl4c38VGPBRe2GckdGWSHx4tSypx4nTQC7LpLGmvHZ/nh8gWbPGvdWugr
tnKBCb06jyQPos2I5vPgz0+XZHKeXawurrPI/EMyj+BWiWCA6PV736gHrHaRPMq4FNUxRxoCb43m
eYYjoSKC/JREMs/LIpHOR/2qu6mcp3O4hA7QVVQIZOsxDIqzo5RPJpN6TSsSqcEIAvc55yQ9unyX
xWHV/3o9yVCtZzGq+LAGiieZFfN6BN3uxnpgK98ZZC7YF4+B9UM4s7fykSOmFEXVfaPmsXBWKMYU
0lDeORHqpQIWYbAFzi3FzBY0T+BOUyw0UA+DQwQCe91TMxymhrJrUfpQOtSTcr9mqAdsDt/Qk2wW
37j91Xusz1r2zxWRSQEHwG/Tdf2Z/MF+uOUwnaW47zreg3Dd6vSXes33qtkTw8XskCDIvsUhOGhF
OvY8G742svg72Wem3Hk1gdm3BpDSVJvffUl0ljL6j4GMFMHYTlfhTHVYFXZeTgin82trhRnvmJEz
wFSSiJU4W2Q+CvtaDw78vASMtppUgpABNalyXqqUC6fvB0cqPh59CcskyukZaMRkN1pw8CPLqQOB
HUbX5rA+paUqGtH6h5Ymwa8KDo1YbzMIuUb5TDHio5JgWIBUxBmwum9GMWPzocUoaA23vtiecYW/
Tf3pnP2GgWL5MeLwXPJOtmZs0RJKFsETqeIw22NMp9tiGPHT06LSMTORhXPUr+EjPVn/S31Dt1Uh
U5zQhXlkZp7NurXS3YTwp46uIcBO8LahD/LRUU95fat/xjci6JNg5M3COmyq7UGa9fkMf6EIsYAp
EA+vuHQwPSusxgnz3xrvwfU3EEO3U9zD64IUBiO5NFFzE+H4dUnCcaZklsn3f0A/URum2m/OBPfq
O06FajK0Fl4xy4yN2gHfv8nknGB2XwN0G+EgDpZtGRFuW3vynxb/lwlTLRn+ebsH0af6sOkOVy6n
S6A4oYnXqdTA/cUyoTzgKzoebEaSYkmF/vGiX1fzj2Dw4Cn1ZsNV8CBeZ0t24ZMJs79VKt3i96M0
iReayHn2X1Y6Xw5ATelDKAYUV6s4FMieYJOYuNknV4wf2ow+vuEyI3DHwPvrcTOx8RyZ3UMBWM/M
Tqq1QLK4Om3JiTveeUpq546JwRlv5mGbNMGb3mxuXJnOAvBk76y6UyaU4Wy5tb/XK4kmMYbMTSvz
yY/VWzPopS3/h5DbS7CzpNso9YwSPCam/SEVOXrFM5vw/cvpwxVwywe2dfEgEHsEKhk2yY0dHHrQ
14mI7kuyMbT1GEVdZO6UCmYhDKVmZdUXxby1TGkvsC5xA9fv92c/8FX3nk0exK0OaDC+Rs2gZGvy
7CMxoD12/YdE6OC7G55IQhg0iPrjQSn3uXMafZhFgl5I9pRSyOBrsGobhykTMhq9gJcC/xiUMwzP
EeOH8kiUffF9zvL0YvGknGIc/gyHqcxuzCqCh5nS8JPOM36JqB41ILc+XOuMP5TnxRblystGYVL+
+MsMCd5tEvOu9LHj3vDPmN9noiegR57muZuqQe+LQL338j1MhrL2hNSzYRSR1gD1oUS+mETtXPKY
Nx0uswAlz4euceonvAPxkh09FAVurtkpH8iwFoYgYOGREN4IVOvun/yBLi0t03p3nawEUfWAKcrp
y8MwdusYrRZhe/+TAHobCXDF3eMw+N9ffvXMd8RVx3A/KXYrarjt4Sjp5uHjvNOX+2vRV+4LxYAY
GjAQokV5fOkFEYB5wbSodCYhuV6I/Jtx2WMofqhzfZltxiH+m+v1auGfWNV6u0xdn6Zpy2ODod+M
yiU4szVb2DH7IPzqQqRwtcEJcdsocPYuQfoh6v8Pt9vjBRf+vsK1FKuLzdyx0ukoOs+c7rIJz3g0
UcxEmBhufvnbqAr1uZAvHPBwRZ4rxhoz5/XreN/EiozK4DUeEumrYBEYfRDn+Z7uc/IUFzqoSspA
R/ZX7AqMXdHo0vIbMF/eYbX5My/wQWncgSzmjR8aZPc++5CVpP8Z2X5ezZnZUh3NoeLbnXgNGW3D
y4gb3zoD0o7RexbxQWB8439KnYTTLcOwkq0ub9vk4gcD8XOynHFMR/L62lpU+FQoQKVTSGCwDWK1
ebcU7HkhGybHXNS8V7CzDBOnI7iTf8YW3RkQWqmmJ4XhCLpwdJWjTzP67d9ZkyyWaiEgMTb1Ty+i
5MvrKq4rTUTgRigES259UG64Wi/uPx8T2NHNRyH0rCkwdcUlKrgcwIfWIEmCegfahkNo6D69XC0G
K64vKwxM8bk3T6RTPwSkMKXfcw5dGcfqga4LKJFA+AEf42wb6qcIiU1ma7+WW8j0K984DBM4NrMG
z3NpRo7aO5QehGMzowGSJ/hJ1m5Ua5lijy5JBkbtRBoQ5XrglC/VjfltOrSMIkk8FH1uvDa4mdaM
7iY9iCPgeNNlk0XFf9iIDbIxBYtzF4bZdXMLcvr8XrA0jGA9W/TTUVbtlnsgAT1ETnOdbWpz/Tka
s/9GqGKriiKR919QNSSL6wmWmJ3qbEbBnnX+AFrPRRBeTtnpXmwIg3W0RefHEUz4Qv9eaaWnsAMW
kLRNrucM5cG1+JG3/SCJ10XXbXabI2Nm83ukhiITlqcwx8tJa2i1tWp6N3QqwNSWTKmtmPvcAZ6a
0KiSfy6yez4ja6UW0eBQcNOjZ7vG4Ee4OZsA4ucpIH8L7eFeeAMHEKomKViVY6AZvdbZBnOb5Kez
/HuEHdOwVUdQMwSLmjHf2C5MycOb2X+Arzm66P83Qx8jb8wEq0cGy5pTdVFT7SgcmFk4ODMrZHJ1
aQ/RK9YLPzPYvwMAXqahSeudiBJ8zFwpxDNYpaBP1q8qDAJ59g58Nwz7hrf0XOR7DP1pA7BEvypH
zDLGPG3nKO+QcG9oVWQNQTTsNz9m7bbkOi6XwgD45dk77LoP0aATAzp+3wKF49uoJAYnvmJGdGzm
FsJJ/PaKzuIbbWdy4k+FeCx5rThYaNusuC8NyxsRLQXvn9QLzfg3LvNS+R3c4VkP6CiYgJCkshIG
WhMNB5UEqeRLfD2CEHf1NA7jiQYZtigV5JGuEmXk/8LSFQjdSTyirE+PRpn3YuvBkt8TMzM2ODYu
W2pM7VRdUYlUa3Bdu1kprTKQXgJ9PMeb9ln1YJHlv2rqIkmZA+aL26xDnLiNYwAHwhjr02A/DtRD
kg2d+JRjFQ4TIlBAS62QToT1TwL64wZ0q97HSE4TP6M9ufinfTMlP7uhMmWIorGyZGYxShktGRLC
xWWokCkr9IxQNkaUhb4G8EjVP13jkx7XWJVW9tHiy2u44K7lbkOeHnSq+tfqXQjaSvmPWS/3Pcog
27JQqP6l3r9UX2yFYPKgPyfmLUBiG1UWPa+9bRI0E8lyaI7Oxbn343/isDqPsAcbUDLyrKfBbrjQ
cd0+CmWosiJB5oxSygQXKH6UgW37/A4Vjv9qpsFPKSl9E34qJB8uWKjnWy53spOq3EE40hXDxEuM
bk0BVVg8ni+LBpB/oi5DfkxVI5OiD76Kr7KGQxohRY0n1m5czdZiq5dqW972O/dq09usRdqWvpvm
GcGMnOleY6Thi9Zfz8UVu6qNbU+fL3B3aNlgsKNVrDRu0LKhJvCigdXPg0KNCsoRNUNTPxxQi4eg
qIOZy1mtwODdkq4oJBZoGMofFISLi0ZV5E7qqRscp3BM23D/YitimPzSsKYUdQbrKpzha+VLoKmK
VQGSbkArSTV19/UKoqC+RmQos5sWWs5bUTVjU5pjP9vDGK9WXveKlpXfmA77b2kTmn+KoEetbbeG
O+FKftPURqO1n19ERqK6NTNyC2Ju4btsBrxZ/Z8oVIPT2i0kYn4piau/glKNklu80NI8vt59QyfA
SiFVknyWY7iMz5FurbSo6SnDULqbDUHPBrKzHAkbng4Bh4oNiLVqx9ytYhJxJBNxAp6Z/CQ7nZg5
WDIJrV9Hc8g6jSJDVVFT7VI7tl/oaS+gHSB52pKlMkUjL5fKovOZmo3n2hddEPoXpJED6f6Yucfq
YgYx8d4OEl4Qe1EaTsfhB5z5KvSSfQeJtWP+otOw/pr5VhY9aov32idLmsdrnvB45Qc8b/h8fFFa
7mV9yDEqyrNJaNf0CWq+WqeKXwe1ceO4UiAaxmPxGWOkggyzAQyhHm752zctgTW2yG/Jz3puutsE
TsoWl5EeSLfLd00D4Bgbf2OHvPzpvsFIUVPOA6FaLJkRl9JMafEORxalOLE0114J799X6Pv6aCKG
GuifG1rAIMgFa/fQYMNp9GR+f3wA4qATWup7PXZKAyidSAutZ+l7XHukbbdgORQKbYWHCW5532dS
R2PHgvZl/JEnSVWAwksnRbp3UEq+AL9v4ep2fGvQUogi9Z88VGOox4NaUDYgSzGQOEriCtbx00FE
oMDi1WZ8TFclZICoaS1j/TTLQD5Rzd96VGzeYbWlmkxdLKGWSZdx6Yubym3hDShdEeAwbkiXsHoU
5a1cHxa9PFVeE6KyMDFcMIMVqlkdZNm3Z61Qlef6bpJblOdkod4HQ3StHNkHoBwcsyHhbUddhKmx
e1wSChrBqhP+GKDgAqWTp1j/xJdHn8rZUr5ymOzfsI5YAa0gW4y9kqN6OL430KeYfchf228N24GW
nwBTupAuuAaD0m8V0Ifzo9KKe3H1/PdRhAcpzF4jNJn41xkpypgu4Tu76CQ9J/2g0qH7ImJEcYCZ
Y8pewf4crG3HXuszxgB87hd8vnDy1GFPgqFjI6SVFLzPDU0WQtOYueyhJGlDW12jnO9oJ7L3RSJx
AUHYfhP/ZtO54B2F0X28fes4VQNdMEiojfxJ7h7BQQ9VZMACuTx6z8pzVIWoXL0xzkPSwq6YbOO/
ydi5+dgttfJAvKYk16PBR4vhZOXWO3zJDil6ujBh93i8ok8wq9z/Q7TFs8X3D0evFCReBPvQIl6Q
m9d4QT3KS/qqgFGjYy45t7RJbKn2S+NZ1IDkuvVbwTmowCCNQGMP03ve2oRFvldsGcOZVGE2s0U1
h0I+6Mv6nlTBf00XpwyOqS6e8QG7SskUVmhkAoz/Oj2kZAX8n6GSCXl/varyD7H2932uLVuVrTgu
Q9bjL+HpUp+mgKEdPLYQ1V4s6yBWG1T7PJ/GITsCsZfBfN1zP4p2+cM5xLNv1ZM16NtqFj/V+h85
fp3VEHOk+wGstE5H5p4SQfVK+YNbKHNKhEtBtsFxX3/SKKiZzyVZQNNO3cPd9lDv7EmAe+ftiYmc
rtQoewgqtq/NRdCwNfxovOPxJyCfFCYiZkX66Ao9V8Qe5tGtEjSN13ZzBZfQ74ASbRA4c+TRny1T
GumTh9x9HtSTt4HF5GaTUoZU1QdsDTkClQKrRF4ZFaPzzPVgJ3WsqyeuUcU2fi57kuQL1+EO1v1J
Tgy4yM0OKUIF5OyjXp3yit9BzPfIVbSU4ZTXEMWwUg+4DNV019akGxBbf51qJMgymtPNXvpci4B1
5Qv9x5jrrK2V77zuxSaVYscvEy7QcDkrUq30s9TqQObUYS3lbuq49/z+ZjHtO6bxIH/VA9OMPcE9
CLQ/YUTM/R63W54a3HUFwca8WpaaWnfr/cQAP3yCaqpbvsNe5zMzp/+JTA1SXprLXmwJjLVLTafK
1HGIUfZ0Du/BIpiivY+MfxIqs8rH7vgnlUlyEv502ovThqMCDAkiyDycIHI4Xb53/IKpsTfihKFZ
f81gt1e6kQ7gGOPZrNVYq8rZXq9NBvw3l3W90H67U/oRWhvN7K6X8e4h8DGcjhhwDSQEygvn6/qZ
YLd/uP/kKKIDJ8zWvLLg76q9dAXI/nZwTCIQg6E+wyLKpNuLkvA9FFd6EbQfcxDgwg19r7Qgzd8L
dIAdHSy2IdYr6iitTy4gNM/+sR9BjTafUt0ATdkVcQ7IBBKrVmVyWC5rNniAjdGU2Clz3yIv0M/6
Cyyqqi7ODV/cbPU9zext6wCGErZ6ucEQ3RIkEmoicznOnvwmqneR4+gAEY6XV0iGzVxsSdhKJdpH
hQccNk5CjTOFtZaqG4ktxHjKin8StSwrH8mAItMo/uK+dGL71kZrE3a+qpJXLoS+iu1ol7xngc7c
hz4bRWVnGGhyM0uZ7MUVQYDZc2l5Ichsnp4+uO6dbQYLlkUlSd/abGOIjvd5Z+F4LLtZzleGeNGL
NHtVI08Y+iLBxlgvoT710z2MFOOyfPv1HF3B8FMlAWZgvP62dQx9QX2+ZjzT16Tv6hwYPQ3C7Np3
s5pgOJyWqnZpcklcErkowYsQwMyV/uzuAv2w1AGnCgf5k+b0f4I7iWPOhRNh7K8PNM+51HkdZxba
6Cu52uRfYwKubOll7WkcvERORk3t27DTlyS1srOP+onWI5kAGjAcPBvBArpU3X4fpzS8/y98FgEf
uOJ2G7Da01CVUhxBukasPlZ2cuYzAVXO0NaXQlSTCA3Kg5PDvAJJSCaxm5RtVE0W1uu/vV/vp9lW
WQiaoMNgSrpgv8CM1djJXU+zvO9x1voIqnb+rQ5VnsNwkkSYxm6XJ22va0Mq22+z01+byWwthHXr
8VMSl7BN+iuHwL4r6SKRY4KlS1ohxkbybIubJnDqKfAyXKgQd2jKxP7ZA0qDRAks6TUAnFwGZm4m
4ZK1l16PbUjFVaNtHlvOc9LfbCdIGxYqCyZhoTL8pDc6KG1c01niF/zsl6GmSgDHml1KBJ0/oUtj
4JD1UFQ6/ohY57YA6z19aqx0RmaEA7709FG3ksiI8VfTyc/h7G6VjebCg3TXM0G4T7hF2jooPqQw
APrHluX1VACJ4L9oHomH6tLg+9j+AQsl5PnX5Nez5hVaGtknJNvrzCdRwrwfYwKO6zaNa3n4kYLq
e6+6qis9TF7c6ye3NAbFqORxiOdYtPwcm0suNTkiBOs26yJqhLSIW3QptdhRYpiSZf1BJu3dX1z+
Mn+GQaTpYCk0HBPMtOPZxp+FTHFJriBFJlUmKpDFXXHpmErnh60L0n9AmCmPa7eANQeRmUNsmIme
312NYrYnoJZTSaP5j2DuOMFjPDa/SPwFC/2umsoD/YFN/Cq72ISK10yjLofq+LMkG881UumT6ecS
iayMWbOfyWkrAF09TZsR6roe3IDgZStg09buMcKDmQ8p/dEAsciin7L4kdIxrK802JBRPXXLHvN0
CJgBGhe8uJWrkuUSf2H7Ds9ojNXrZiAnseg460hJyziJz+iX/sLJuXgagkKQFhmBlgm/7ha4Gf7M
6362zXJWJlS6gLvGGQNgHjBiLtIqsn40iD6bxO3XltqZZxDMlfkhdH7dQkw932j2+6YiQazVje4+
r3vFBhNDXMCdRNr9xKnR/3XbLVDlwtG3D6INy7mDf/MJkHv8bPeVN9vMNz63Q4vPErY2oNgMMWdL
CsWZKrgqDZrHef9lJnV9KcTJ8vMrrcf8lF+1gEluD2FyX6twEOTPb6sG43w2vxj1zr49gZPEcqtt
bFqHbZwFny5ElZXJSrIBLxzHcUATZ71Sh53rbrm2nFDg/bDmb1LAgM6LSeid3LWhu2vMDwxEuSKt
5B6zP/GlRUKY0Ag7FEevtZLlqPGgUVg1biAuMSFeeLNyxAu0HWJMHVZjCzqIA9FlmzbP3z1YyduY
iLAtoAI0pqTmVv90gza2fLiSsEtvFQEmriuL9e33X4Qnm8TGVMKOwg+lctu2e9nLpSr/E/lI5MDJ
TksuMml7HI/6pMonbCD06FASw2LTfTIb1Cn+LYSdNzp+RemAm9xV4xKW0VkwPOOZZSoGohA2X8u4
Uuc9KhhtR2G930Xog5TSBku5Cmtq4A3ogSy2ppeJrJJD/Hn16Rbn6gT34TaLHrihQ4MChK5sOKyU
wcMoq94DiOCuKG9nWpsX21YNQZDdlxcuH+PIF95EvjvdmX0wcTeoe9afl92UlUuhwl1WdIkkAOtZ
W5V2n4TYkRIAuF9DFQ7w8elDyDnouvDgRyo1BhMaTKPu+AEJbwOZXZj7Me2w/JP91a1xWT6PzZ4t
NTwabXkM/JZDwVVLrnI+Rme8FqMAybgX+9v+nHQ0BiZYvF9vItrUKU5jhbOmv6d1uNeqL8U48TTJ
KOinhsimP5lA9sxJCcRbHh/IOp4tVGQKQ8ANnky0ydh0hJUrndaI8JqvVa7aDlwQaHMQWpkEU6I/
YYsfAgbjGT68hKo7sT5XKcJ4rc+OgMJQNw4K/36BxBUf+A5S6LjwvP4p+VE83Ag0jJYIRN9S7WE4
g+3seT2+LXmxqnEiAloxOoYhVKy0zQXTlCcWfg7bfFBxxtDh1BkMo2Rkxn4SvV+zrzDe+oGa4C1Y
aEMKOJ23cdNYCO8CMYHeZEcfrYGc2jKN3JtXh63N9wTsYRmQQ96zysYytrqLomGk+SNuYDwSHQcD
1jqlgVKf43fGfJHRO7qO8Ip5TSBE4TEKgJl+caDY1iqxN3ej5FozZP9LLra42D7nAnW+66Gd9REy
MlgLKTSiwTdqRugoFrqJ0iBCXD5vVTzpjEyq1O4lRWTgmwOpEBPGSLx/3vQl0nvU4+/ve+61i44l
KIwXnCx6p7lOMXwlyoYlXal52R4+7ypUVdV6LX2xKG5D1aVPFX1t8rz2rNEJfaPfZsOZP9MfndB8
RdtOdR8BpQJ3nkZ2KSlYnbVKR9S+M+oAf9A/jv7R0s2AYVLQryE2ekCeYIrggJ5V6pu0PshzTLCd
Te+KWqXWbLBZikwwkfV4pI4jv+kEXwq0FIYf8+n2CTTNPsu2xydXVY5X1mZLyvRUCljTafNR0LJ7
ZenTbyzvJA65Afh3KdA/PccAQX9lJYrWsG3ESXte5dv7PwDpta4meGzYHiNmu3C8N3jRbnVX2NE7
xUP8kLI01pUXqQZF0rokvqdL6z1xi6VQnRQxK64GDbiQ4iWIh5B6o+t800u9Q9A5Bp+iEeP7iZ+v
NeQanPeXsF3SLqIXzheWlteWhi/lu+7+iAO+e+HlK3qR1HVaV5KAx/FQrAvLG/3N//oSNAnVqh+z
VnFMk0/DFWRMcG90LlqpijmvMPhKDudtzK85qn14sPeDmCb9WWyoymKjKdiDmMrYXNt/Aks1kLpI
IpasZ862Pr3leazj/DFY1/0gvWWPFBvzwdhZjpJaHGLwBwF1HWUmAALG4rMkqcKxk1kqljCXNyaE
oF+kwWvtTehYVrhoYtK8yzObt/e8Jiv4GimQ8hct0hGUiwVQg3tKeEBIDiN95siNnlx/bZ1iirch
2p2niCrUmuI92VjcuSoiIC7mLPY1blxoeSCtHSyz0D3h+IWeaSUk6QtypZoZ5sZ7HQYCJs7UUM9b
KUiNBIb7UoYGyY3S1xyMCJoZc5nEvDhDYe6xaZ0VJPrSGxLn4ITDAJUcwBTWXDvOYszGsLqLbl61
ID+7Nz2jt6+0qLmB+eFx6iQZ45ThyjErFsykfnqF75xzRWEE9Bn+T0WAbYwKkCRFLPNTqWQ1aNTA
z2nMf/axPT/HnoLwhaTvKZESqPIjB6oYPShSW59XU8S1rA54mrKF5ovLoV+LsO9OpwcohpAZ3iHG
YjVPnnO7BuecupUUKhw1PTl3gU5Gx5hHDMWf3jBb8UIyYtNcmtWP7qUv1KxSFUzay3ClU+ApvzAj
069w6nUs34BUSdKMvHkOGEujFhrTIENhyG5F/jwi2tPN2ntJhs3qtQdNG4CO5b9BU0L6bdapvIiY
o3qz87MJTGE+p06lhfLZAaOiKu5XN83OTnpXENQZH5hjVct+bKQFt3rJE6YvfTuPzqYI0KnhCrZZ
LeLkM7ceXsJuGYqHjVIJ3jLR2bTpuX/EE21HZbTw4UqdIKssC8aL2X2754y8Xj6KXxgyYP5Ukv46
kmGLmbNwFr9P1wR2VXrBp6Voz9PRNFddszt8pR/CjN3L57R8TNOnehelfIr0JxdkOENb6oEnoulN
K444Guow0A0rzqqkoNoNkWWrPS88Fw0XxRS14F9TuKM13+y018qoyMeBnZJRGFnb5v0gmTkmd1eP
fGgs+oEUxo5zzezCsuIQQh6roqMrt+LofqB7870ID3HhLEx9sk7iW+zd9e6kPg15H+MV8TeKQO1z
UaOIyC2GB6aa4rig0fjVXWoA1u3DzuWrFPK8czS7Sa3Yqd0vZ2gwFpikHsyD830iigGktjs9EUxv
qhL/N3uJ5C+BfCP7hb0ll7DTvqJcRISBWA3YiAnGcHobSkaUIRCXPm9kxX33B5eDtnI1c+4jc4+k
EClH381M7eOvBGUMV/+LDGQoetlU6E/OAnLCQIBWXsqNoNZ3OFfm4WHeHnVSlBr4EkDgQP2P0CMZ
U1oY6cfWOFzo9U53I4goYjlqgSpyc4JFfWyeGEs6Po0/VF8fyN44cyIPjwYTQQajXjneyFZ5yFQq
QLUXYmMcwcmyhcGS5kcX7lQx056o3Jo3PdsrZfo4E7IuuuYGNasTcqiCqwzujCFW0Qk0q/F5ly7C
mAPBktpNpiu03hGEucEQRxxTTtcmMKp2rFFEpIpryF8JsVP6Dv08Iatr9T6ssVWYcVR1tSbqgfAF
Ax42yi3Jfa9YAnp/lmE8MbQgfMYVffTJx3NlcAsjPX1atRS5VTFbcnmMwH8MWp3skVtnMjZm+sdm
IzZGNctp3Umr6BYwwpFSt35rImLw7T6Ie5CODj/C0Y3N265YWol32s/+VSnIXaHy+jJQLAB5d4Yj
2i6oE7S/w3ovhx5cn1Biuyy/mKNVAgpQwvmWyFz/FHBJruOGljM47xv79xC/9DzaFjts7fSrFTh3
9E+wkNpUsbsRyDqLCHi908Vez7mz1YxBt8yuBUrYI+YjK0Q1Qht2agBR0G38jD5oI3Zs5TNxVyqv
+cP7VyxndOhPj8jiiQXzkAvNDQBComTIf5S86nE12w/Fk6oLx7eh8ec8g4Qzz4VXtq9i10F/ipII
suS5VI+lF1Fww9mtUKsxGDBEuWgiNpp/VfdroXAzyZFlYSKKzta8IN7p0eZrxViwTQhbSlJ/A65R
0Z4cw2QyT2yXwJp54DAmBfrxpULs+U5uG4/UzCs5m8O/PYUg8zel6pfOETVMycudx8k+ugQsZvDA
ZCHQx0Oo4zvzsXLzp0VEpHT0kQIhDuIvxUu7+47nN5S2Fqd9ijGoE0NLYALOGLGxuZAH/eEy5HKp
RALuqHZOmPsCwdHI37QKJWkWvQbsWhN2bPWyP6alB+/tsPcw8jYShk52j1Vve+sW88782g4jyXyl
wniAa9PX76FJkPvhC7IO0HpoEsRVSEVNpOjO38Y46EX0oQt6JH/B4NjWJQBhYeWf8Zjr2SROjxai
dBoUDl0WGWNqMiszgyhgMIj9SYEyacLlb+shbnHIi9GC9wheKFCoP6rkvLcRUjwL3GK8v2ehdIHI
3agRJ3v+KQr7maMf3JJzq8TpY2xO3PFfnQtXWEPatkIrW6okdFvJ3+WIhQKHs+C6V0EkcfcMfE5y
JeOUwSJDDSjOr8IqJ7c8vHWlo8hlrDSeNClJEeXLSJ8NrfhaomI91aUz0JMP7ifWWK0u7CTEXi7V
vEfFmi2hTCumL09dkQOmaSjNTUeeYAgrH3EyCWzL5WCWDJtNswwj5B4i1WvjDO3O323U/MCEtAu5
+SlSflro/yPYV77VmL5724aJVW6EeYMf8QbUj0pxT1hzj/yR6Beq1DMPlKSp/lschT8NDMbRNOzI
rwO2NcZdx+lZst1SYAId5iheEYUAGFL4w/KegmuU7CA8E7eKy6/uS/pWhpU4Ytpk2cBkaHgSEQjA
0nzEI+4iAS3sdk1inDDOS4lw490dnshUI9aGcRa9ylYSCLiHxJPAY1t8M7h0XUmlN7q/K4XActvs
NkJ3pbCpw+onW9l5cK2d83ywuL2Ut7noZER4ZfYnEdpDGyRbp5uhWyHtudvt7pBIlK0dXq1pyCVG
CpOTZfLEuSi99GxWU4S5n09odXQ+Ok7ZbTKUBhBlxA+R81y9X/mcub7XuKFuSu6nUrRonjC7r91F
FC06EiBA3slRd8Hid5PorsIAUrQ1lxWXuWYkU4CSVXDFvCyy2f9JDpgxSugfE4JVGk92RvV7euQX
7lsjx4JBZMp5RBuNMoDYl7C79xmHy6lpAsjfbVU9x60RtryoDsNsCxWVRoJtk6GH4Inr5Spp91/M
UnsrLPTBKqmKhOUniUcsm+db4Q1R07GeZAlUXHUb7famtSWoFqP7m/+4mwflI3dPTRtLV5e79qdo
kuuvNgSfBBQYZFYbHUB4AEkrTYkVMmvGPmjViUllXpaVrEjtrtRhUMp5pSN5YO6Op1C7O6hkhE/P
uap/rlo6CdUd6XJTB8IH63PhlfwbkO1KVY6vV041WCU3tV9Pfo9SpDAjuZvmZWd9cXA6iwjGUtik
nAbeF/3esETbHCs8to916EUSIEUl5lWyXfWdQx+iCccB3gWodgOAvRDC1tgQT1eOiZ2l1bWtOBP4
97lxqlNmw5J4yXYgHXptwvbF18BSWT9te8AOU4i75ZE3RwUrFx8VnY6yIczeL3ZcWQF2Xu8IUZai
9b2tRNAjPk5zwoeS7ruB9sQwzvDyFjv0b+x4j+Vx6APW7Jx5pGdl0GhGBkyu/iYhlPuJJji1dAU4
upRmgAFrrtL3xfxxjSVtLy/eRIISCI64EcmlyXPGYG1eeWthQ+xDfPv9jIOoWKeRVN+1tvoUe3vW
dnFjl/WcaB3DRpy9yc/H6wXRraCi9ZsMvZfClIA1f4fztHTW9pLc0i+QRDVr2isgji31NOpWmM1P
9xvCaPhC2fjLYe/PwoaZLg+pUIwTNQhxYYVI7d8fQnofN2M1bu/PJrW6aPhds+GlWGsVaDC0aAH+
lX0rt9EdHNecIVVo7IneNtNP3fSAeO2pHSzKXaKVkpcnJOo47fHACsZ5y04HL9PKKqtb2fyJAVVH
TwUSZl/BPlRqa3iDZf9UPzPbyzYUd8efbNzEm3kneL0T/J8b1Ye09S056AiZGLtNwE/pNwK6Dr8G
9euB8zSvyEN5Q5Rq63q0DR0hL143V4af6q7i0QCW2zuT5ADQ4oR4MFAoOSvvOaeVb3gWAXB8aZcF
IEXM2fJGtGdRNgoJmeAYk7X/EsMS02rzmw+T1MuopUyOSzY5Cip5MSrl860I1GxO62PEL4dsIkra
fglGuyoRjpHeOgbrxhvKuCk+Nzib4A8VyyvhfZsH4nnHj+MOAiEI2vG7fpxfPpKyieC+nReW9pOB
DJrQcdJ+5fXgNXulobqlPcU4hwEj7wmRyKxYc9osAUQGGd3Zjl4zLonqTZIP9DPJ37eLi5M6qPKI
JV4yjLJ7eFL3i5FJ0cebiJrfsZ7l5YjoWDhAsCO+i3PfarsoSvwN8LUem2jh5D8+5ArdTdtLnqD+
a+6LRPw+PXWHf53NktYK/uN4zHye1TCteKyajoCVoqHWUDB+tzgFk+USorvWvpHG4KirV+vsxAx0
YX+B3cy6JhS1AOzHUZGLfln9QqUrEbdOocc7SPizmbxJc0EJyMW4WmjFctB6ZsW0MtIJ0HF8PMNR
m9VyxcqpxMrIHNaasL8e6t0QylsC8X6IKkg/TLfhY0YXiLaDyiERrxgWH/kQmtthOrTqIcKntIZA
mD/uLrs1FNtA1Gs9/Xzr4kp9FFGxq7ywmRKrZ1v8bmhWSZdeO52r2kizN1LSSjywBpLwvcFCeKP7
QrY3XkmIlQ1XMr+v92hDc1fMfFkeW7pPjqmX51mZglZz1JtStYBwHhxYTtRbMhXyMHSPNXc0/kGr
GmcwrRPpwJNVnihD+k8Sv89W6QFPzICOYtsKWvRRcpgf5pbb6ybItZcSz5O8N5po7PgrD35OO/7A
1K8DYw8kIl5L42lUcjhTZxjs8dAMxWuyefbT+e6jIv87Fz96s4qpALh7MeZgce4AUQe7LuXQs0Kc
LQnRhOabGJ6LBwG3NffRzo2PevpmxVozufBw5JK7DKwtvHcjT6Z1IIixGAgs5CwjbPGSAQlItCcy
KNsocfkBqRaCmKeA0hIBN3aGHY05UlZraxzLaeG2BIHw31YwhCZX89kmhpdtXo3Eup2keCNHeF00
8onMm95n7jMaIIxrPGffXeHYGnyTcsI+t1QV3GezGL42JJmQd9yCmNfqGcLAeJeduKd5Ums5T+i+
8ntqFAY19FiHIX+lBGN3Q+u6JrXFAZH6p0HqeLwOLTBdZ4NM4kqLSHgJL3E+GvVOcgQtR7hzK5Hh
HPWBp8jtrUXxT2WmG4/E/NU3b3nQaFwXuhW07hde80Mxjt8UrOti26YHZPhedjfHbQixGVwuDKR9
/pv0VNLsnWz0v1NSjQQZMLPwkiGDiejfrztPtOGDz+5ssoSFGQZkCOMGZxlbeWFmmaC0Iw6SEEZa
rXwh0Y/SbzGl+O4+hc5cnT9wRPYRt0Kw3P/lYRJTHtN6/hJAT2pv05zzvcj0WSeayjQrOC7zPIbN
BzoyTgYD8u0xp9y6MtpWmdbPzyoCwhoGs6AVaalpWaPTqgMrGgOLlns7K+xJegcRpVvqB/Ptd9Gt
SGQ878+4SeIWtWhUCsCC+uTlZe72ie8GXRPJTlgVv6XDM6OzNTuQE1omGU5Xyi2KDqKasbAvRP5D
XzT1cLMU9DCoahNxq76cD4KZ4KskNkoI65upHftalaiBK2ix7Gh4t7Hx9yPlzsl6XdrtSDjlk+IV
qvBpjNf/yRfdHaa6MYC3bYCDAfamuokMVnVYjGKLl1BvnUvk9WxKgMe0JBI1rZS9fFaE5OUnZ4ut
YSQ+7fZmCxoCOIedDJ8tDoCCFuc+CmAv9vReFCmKRquR9ositQNMQwQTzvabpaYVSc/0ahOnCXQ/
ls++Ip3vP5CxdCs4m2ilOn56FONICL8Pq/KR2m5hwexnhvBZb1HYkDt6SxYmLW6rQUtx7IIuG/EJ
PzY0QoHdwi377l3o4YeXcKr+H5IMOvSJxA9USQWBhpUZf6compQhjXew8zBi2CwaWRp5X3lPYAsK
mbMI7skbkaCkoWiivvzMbFzQiftwtlxPlNKQuyb3nHxCz48GK3EbLp3iCtMX0k0HXOyL2CfJmfhM
aceNgc+9DAn+tkL9f2Gv8sM/onZQ4ApdGWY6ok9XwiQs+eTehlojBiu2zEY9CKYER44vFG/8bVJg
gwOp/hdRR+5yfpindMR6556bjaOwk0it/ahhI4gosBLE5Er7J9gqKXTsN0LEzGRHGRvqD3y1wLCZ
B40tFWWBvrxceeNlWOlJCbM4JM4ZYv1kCRuDHSCJrUnDuuW0GogA0kvtULSB1saDS9apQ5j+OhKg
Kj+DeblaTh8Mz/BtxZeJ61VHBN0Una89ixE6B+2OaGPULfkpnA3DR8VSc8PZPnzMee6LNQyudSJ7
LigJ0AssgjI08gIgwBheM2+2SHQAADPMmLPFfX9uWJk3cG92MPeCAZ1J/o3wv+TlEsJfj+bNrNWN
0KdeWkcyPsfg1MhWe20r/00OruSNb5PQvbAF1BHGGJAJ8UiCaiwKcEsOURiqLbs7MPqVXSja7G16
beXtcBWcdotI9Tc0UvMaxIg9UP/FVSVxS/l2k3nZBkYC431S8cnXfz/dodY/5M6Wq9dh21V+Ya5p
ytcjiLWuNclFAoj2Ea14vKt4j1SOPgV7t4JR3zmCXEbUQRE43kTRhXWUHZhc6gQryXVSeiiD/cEV
1Q783D4/vm3Xk91Y10wVvsFunPK+5JCcH7d/Gh6pEAjB52ZIgZSW1PoPdfo4bqwvwTzdnkKICNLN
KWYTYSAd6SDXuqus+YjcY+mgSKxjXFVhYeeky5fK6KsYOi//nkhuRNoZhd4W7MuFf10s6pW5Vc66
8XYDhoxdQYFKe8BylaYql9iDFeSZ8F1c1mRb61oyOo4OWBfsQfNw54cpSgIAIahI9dnsCAH5MrAT
5bWvlZ4FCnjFlN7YuF5xfLT4IaJDHvWBMe2iESa9EhwKbYKQR9ktNADmpI4Ve8+LLRopXI9SMHux
jdYMVhyRLr4exHJTUhtbqGdh6e7dXNyQO9AAhgCdXIm6os9JM0NN4JKZ3/GT6DsRrpbnNdgS+DeJ
4Wa9DFCWN0d8P1w8uYQnxKZXslZ+u32kEF5gewzfKlm6CQnzwDStkBwF6uImR7wWhBfJNTPWg5Ir
6XOdk8odkgKekwpLRaii2ZVTNcqSyacXLRbIMP5p2IBZzLIuE/ShJNeAO8OKe9U0x5DaVz6XqsNT
fofrMpOWe1bhzkIhok4aGLQ8gyAPgSkSI/v5L9Zjy1NuIbUMAJwsm1d4bwutLTeH9UwdP2AfgTMj
S/crgTzuRs0xcEGMGMjRmkACYUfDUa6WJv7nx4iHFVMTcViq8pi78jg8DFcqPAMitfCsMTUADc+n
oqJB57OGN/8GQepvjTpUj5NHcHpEzZZCieahZGw/FmcJ+3T3BFVbBzadD2dCooNAdfhHBZAoC6T/
eW5qB7V/2/g0OZFG+6fh7Hy2+gsnvoSNnQexh5C/WlUgAAQxFnoOHpZgiGlCP8g2r+VKaSB3+L+7
4GSzEK5yBMggmgFTZs75422fV65XnApf9GPlNLuUQ+TngmgVx0gQ9vykjHzpCSbaWwREnSlXPLwC
xR9deDsgOMmKNm2otk6EPUDRmULa3UmYfiunVaA0ainDqZB7d/bqfWc8sKQcGGecr/kZE/6OS4WY
YhZBdhvxO5bNdastfnPaibzu/QZu41m4mCxVVZRU1qJK1ND67BrbLa63B2FkhDkY2s7Gas3w3Sbb
VM3ekjzgRtk0yKbFO9Ney0GBDoTJpPGd0D17BVYRpH7M0ROXkMO5ZKr5uom6Cp9hSP/VMuShjXju
HgtRD+wfm9Kw6+nfksr3cpH9nzbPadHfVYejmjEzl6h5SDHI7Awqq1vGndCQwKY/Vxily0tARvp9
LEIPZHrWuVWcWsyMrhokWJdlemHmVO0Tuk1Iwo48fQNNozbEY7Tc9WbqBjVCFlt8stSgQvU1ijRd
4W0/GLR0+tcv6aGRf5zE2gCUiKO31as3aNm9r+wPOLIAjESYWCT78BU0RZT/jkDUCJs+b7/nCCHb
+yJGTWNwM1RbQdQ+T3Pb61OdG8lVTxlbUys7aXZxo8kJxDqkhcrY/91l/zK2MQFUYEup0ZpsbUGT
F15qcBlsO6LRzgd2z/z83VaUDvvDY3h70L+/U1UAdogdjp26cO0n7/NwlhRxYsmtXidkCqU7Xa6e
FldApBNtp0MtP/iPpKlK9J5u8upt+/r5DqOBEbXPhjjMdtlb0pG/eY4Q4rGttbRl3D2+VAzjgL2U
SOVu3XMlLZDJ63I7Uavsxytl3Sygq6bpNvxFDFCNZ3DE3WHcVDM7iRlZfxAtnjgxH6Pi9tNRt3uY
SDC6jCHhK2+9Wn57IedR6NH3oCy4PWd8xmKy9HiNzUxvfUcc6nEUiWQv1j0cEy1Tiq2mjk4Wu5o3
v6aPH8oxDONXaxaSKNvsQYcNyfV6emiAXKxL6HHcQ2yrzSEt3S9w+jP9RfxRf/t9Av4y37zpYZ57
TSUsSjhQ+CJ6+Aacrdzx3t6IYLLuGyV7unjav+kRYwxtencevOs/hSoomhxA2mOeCI4xwbUG1CSu
AUZ0wgmgl1fcm/DUdPx2aMJPuKyrvJWUPa51dduFUp/rald4cc+pkdanF1oWcHgvmz6FVIpu+2W5
sLrG36bdGfJbXsL/kYHkshzcc/8JbJ0wvH75gAkvaZtk3cPuZdN6X3gf0Qq/PchkHN1atjznlQx4
Wv74VFKDow3pHMIU12NO/5eNZkp6J23FafJ52dXBGvciaS87yFLkd1X0W85wnHlJR2jRGF3IQyiD
p8YqZhWeYE3Jq+k2/Lq88CFfqhCECToV595/K/Z5dRpoVWJvrbYZFnNLEugp/Qb94t7c6cbFY9iY
DPFm6yUjiFr2lsBBrSPdLNq1Jd1EPNtBIaN9egVBQDFmAUQMdt4mYl9WfL2eavMxJTCRAU5Srj8i
qncYAV/3Mo9IXPJ7CGsS045I4y0q+VstlmP/meseUTtaW+FdqPl9aes5H6zqD8inXV2a/UrvG5ZQ
1GoBogF1W0bOJ2zimnNFPUewIxbY+nVMLl/z9I5ZicCQDbmpIjFcx/Ey7IJvaXl84qCQEK/ZMO8t
SsA7ghinqshZ6W7l85V/jAimUfE5D9w1wP9L5O6GC35IlXfASr9wNxnAGBzWHsWMSD5TZO2Q1ro9
gTGxRcq338hXHTt6tTEAbbfuyQ/Kj90J2XDzOQPjNe1OMDcLAWQGOI8H/7HVlihXE3VN2BVlPGxN
SpC/hP3mKNYUxy0evb5pGjP+uGaA54qB1S80BxRRjN0Mfl6N5fMCzuf6lrl6e57DSKQT8dVpWf/w
LplsIuvlvwXy9G9MCu6omFSdWws2mHJ2hPeCrxqrcZu21PaS5kKQNLBA1qIn2KkFlwvCmQ1Lqv1e
SJNCGtaFQLmqeMExnuH7Tj5nJ9oTN+AmWt+HemVikRkUX3+GOjoH9I/GvPlO2D7KKshH1xQ3y8To
8Tsh+Jf918EHAPJzXzM8+Zn6xE2IPq9V4+4HOB0klbJntl+5x7e+Jkae96/60IRp9+R6IBSySdvj
X7VAqSfuuUl6hnh3Rmubq3FSIzdvHowN7RoT8w17b87DdxORzUONVzW5R62anKUH1tvmwTHVpXrv
n5Hapzfb/tGjQBvvurQSd/Icd7I9XKmBiBnZ0tGY1xvsyiAo+DKtuu66O0+CgGeOOHUDCGewF3nC
Ffwt2E6Wd1zggrzKkT/6ObP32pEFGlYaHRpSY34NFBNwEZEVkOyWE4sMDW1Jz37ZWG2BHPALXBQ1
33oyPj6anKUYsBWEl6+k/Lvk37r6WP9OlzRa1drBZmIgoqU5WHUBcX3ATfXjdscMWwhtD5Wqxm0k
kCBbK5twpQw7Y5tTTYTlC7Kzy65CD2lB1I4u38hZxLlfv8EY6NR1yHXRP2+zcQndv/kekgeGfmS2
OZYbAt0fdU4fl9Yczpqgqxo4o7yrsyH2DLMI4YL9ApvLeFbGwJavbHB3Tyrdp+mnZmikZAZhZVzQ
BRln8DVq9oC40MgyiY5uUUqj0FYgTBTGST+nOZFZ8eYqePP36jiE4KTNoWrdQQJ16pg+Qw5eEHcv
3IJy6Dc1WRxKn1CPXDNvpT5Vx5B+HlAqCFhFZzyEXsQpBLSmBusaWy4sAhbjyJwouPfNEHLuCwg9
o7mKTdl4eO6LVqjd/bppRAV6cTHSywyczNSx6xJH0ENp2/tB/Ug7/i948XlPFJEsROMjDpMi4/B9
xp9bR18CYajMEoIoNqD1WVz+vXMYBZ4EqbozU9Yt9bmRoKG5P8253A6JrMhK6g1H7xkKkUU4+QMI
zvn8enyCxKNtPLMYI15g1i7sroKAQDV1gB162uhVKS1VeL5mxSEMmZ2JYyqn/b/kcZEtYCNbc9em
NXthyRV3lL4YJtO4Sl/xyPQTefjBxsWnSl+IKu5AucrjseEvrnLIQyYh03IrLQR5mZuy25MwM2Om
tsGsmXoDalGuhD+66pSgfIW8YK9AeWNnEek8zbqHKDYqextbZTuFLPPkBLLGwNajawpXlyS0ipXJ
F6uKX/+9eVu8qpBXCsCIpzZTTivhVVxM01vvfBjA6T10FK/w4LLPqSfYxDSKdb+w8mgaX4yoPouT
uW/bCuHgZaZBxQ8pWYx3Bdt6hvHjAWyiw4Nbmzw8KU9Ds90ityqOQZ/ZD24mOYcZYAuwxJMCifKm
dttcJbXBalf7UdL+HI/k7B0q49xjFnzelwzuw2aurH8ThVn+kmbNTCF1rjbAQqU7yGAU99roRW1F
/j+SKJ45qHfbQjwthjq5ewAvNm2BLExyeNx0B0o+CsN/3C2H6waBIU3RfjTvpUXMoMc4jRn/2epW
PzVggKkHOxGcKTzf7u54RzLAuHuFxzKdKRCot/0pwq0QvLE5v65jwsI4bEaTjvPrbSp6gy7b2ngV
0/s+ztPaInKuJNW7N/H2POS94mwEJwBT96bUs7dLKfJ4JOonwVNsJYQvxbDz4VTI/fQY6pmIgf6A
SEuNrpMBlOq4GVlx/0qXFNvs1YP5ztoV5+PHBfSzJrTbv0bXcA0xBmNJQHPMNu6/cUKFas2Msn7m
Hmq922kzC/uCmPze8VQRtWAr21HfhV39ahezvj8rXP/U+Z94pYxPrYwT32DpGhb5p9wHsCZg5X4e
+BydhhEnrl/XNUrlsK0lT9taQmRCz7+klrbnwTk5ebu5aXo1S1yn0c9kg3bMy/0ZrzNR9aiqHAeR
Z66NqpUlKTpckNsDybn3oL4FylPjvC++XX8RHMryWc0j821TndAk3F7bdgJsV7djO+SV5B3PWlXh
CKH6o3GtewfIgKsLzmFeXUrntGreCe5iugaBc6/AEUOcRBxtz5frzwRzWniq+Phj1JiElbIgIxEe
y9lPW1jp46ukitaEc2xDxV2k8GIdO97E+tjDiWdcM7mNmf43feekVOnqP7m28CLnX8RbVfFZPXb1
YJhT/E6D4QJvEUuqIvvFpU+8Cx6mGxS08bHrQ6Xp+3TS1Ztj1HQnOJ2g/a36q9/1WyTOWkYfC9wU
N3vdJE7Ffpzm9ROK02pYNDHWKr7hwRZ2oY6Qzj+35ueCWSUOJdo8b70if8ie/YfrtaAAK3RLFlbu
bsXZcaFd4KV4In5ixWrhIuS9/ElUfwZMn6Mn62zOWCyZR58vvQkpmEFLwMo5nbbsxss9xp9vmWDp
pdM6ru1UvSNQPjoMP92iJs4EMntvrj8BbV5MHPn6TyJh7CWC2G0+uqnmyLdWfdN9FOEu1F0LkOf+
2HhFE5aBDh8Q9hIavNWjQivFpvctRPeHyS4Cbpo5BpV7NJd22QSaWGcRuLhNRd0+6+lm71cwu5Dp
b+5qRjZ1qB1/0hvtzZp1S1OAJghfoYgFEpk5cd8hHVSD4KKqB93mnlJUSy1E+cZ0OogZIqvzvMrr
BEs2BrChPOdZjf2JvOXNRhwsP/iHYAVUHzOges93X3OPydMo/W/9QUuvH9TollhLg9i6euQupo32
7FZO/N8RajOELEslF1w4jzu9cB378nSiquDr63ttiWWQAfw4bKl4cvsXNh9DK+23sDads/PfFWWT
izaLKn9RGoVUQRLhW3B1dA/pdQeyAJR+X/Wn40p/H2zSBB+nYTCcFboODMUOo2TkCPARR3T6VY1I
BRlMksKtih61o64AivNnTH+ujOoA0k1QKIMy26wvA3NKMm2/ZSZpSstyXe6Lr5NGQ0a2Kf0OJvwu
j+6zaz6VG8f6gM8CKAwjXkGBElhmn/5eFv88oaKGe80njzRXTwGZV059NirDU2jLz20lqDVOGU0U
lA+reURfgtmXyqzSJK9zAA9lm9Qiqop9FlGxIyy1oB7IOlIJvzzr4/tX5ne9e3B3On+weqF0J7kU
hAhIHEOs5SZ09Vz05KdOPJdgxrkzf6IPVtSaXyacuvj/paTeb8q5wHht42xNlERFQoZqauNWVVQJ
Q05lz0qkdZ+kmRomUIPZ0AAo4qgP8eLTDLSApY93y6NgFEaMCIaikduLHvVu/YxnoI8fCRXwqJ4y
CoX2Zu2KNnjHXha3OAihGqAcMMb+aSkjrTdo2KbJYrFgy5rTxzyoIF5wvz8o8AlrrghsI8TYIqai
6hnOZm9A+9zoRClx28q4dukl3kHN0K8cXOjcwIsNXuZkldgzRrwzrNH9fvkUfY+A6FLpHGGq/8Eq
JhhFBXKCKsWeUL2vfga+29tOPBOatrIuepM0YorEAdoOdn3hUevgZKGvyFOB4zM+2dsohK04c6fh
FemxYaQCiBHum3GqxzjstcReYzxKHt8Eje6JryhRo4F/KDByQZl0ahZjum1IPESLkQck4M3+VBf9
mkXyq5RxTZkYZJRN/C8ySuc+bRyT/3I+ACmUfR0/L3ifY30h0v2rnSi364eZAz7BiGZFScDtMZXI
IssfYA2T/eGLXZS8+lZzos3IgjRuo5OkdxSJVhn7fhkOCryM9t71PWGIsAcJwCJyK2Ji6ZoSVBEt
KTVaNnSFYkowqnfXjhVkThy48XcPAjh9Y1mgheM32F3beV/hW+Q4Z4VK2Umz1IweuEd3Cd6ocmSI
tvxN2G34D+/MfJskfixFSnlAxWM8GxoCBN3OO5E5DXQs9iJ4X/BSdHU5DoP0RY4wCEiu5/9vX1Qs
lVkQI6GiMpngd8YkGkHglJY36I1phCEhzVUw53Sv789rNErt8UwtwK60pWZuZ8cFsgYTGGPtVZ+h
mEVEkYB3TJnhWWStWFxigecLDNh8cedfo04Pa758r9kQwKzxV9ka3xoo8rBFIg40RP9OSW1qBv2r
AFfh+/iyDz0uyHZoJqlv4uZd9Nicma/ovM8wi0TCNMVua3rrQ9471K9SoiwiwdgReeCzPubLJZfR
9eTQPIaPdMID7WgPfRIW9Mpxu1U8H7KkT1iBhvbsnkhCfl2j+yCiLgwl9w9Hy00hmTYq7/hckVZ7
Qod7D3ArmfP/1QaodA4B7U/o/vpdIVXyWVi1xlwYeGtiafhtKXD0JddQ34LXHr0Zb7gcKU/gwhXr
9t5Pz2A5SC3YcwapAnFM7fB82g08tvtI2CllsjBWmTONHjwP/1eSGL+GKNXnXWNhRsY1LBpJWN9z
9JxQuXmjR0OQvnCDnf2WKN6UzbvOKU+9hNGfd00L2fnRtnnOVpWYKE6drNbloU5AHo+ct+DJhFrz
MC6/ObCUxtdv02HxKbLRKHdkbpyjfifsOAqpTPXQsY27RmKBJTkC0VwcBO46jthN5seWwftuy3Ud
tACIpnvQ+IsnyE3DrGOrhwCrAsYOAB6LjT+m/W6vyiPCrAewbraDHlcSwltRH18WmnOwCjLbcYv7
Smkkv1aEQzIz+rYeme6YIUE73Fi+p3uX9CfK81QE4Uvh4uCkGHGiOnkGI6DnpuNhvhSt45OKUh4K
smSjr/i3b8yaynGz54rojejz2RftnozmL3t09e61DI+pGjRosm3rAagNllRL2kgOvvQOtQT2iEba
i4zrMdQDFbmCAMPFBl4oWjI7kF2erc4tT08rnwtjBnXa2JzUmkeWd7zGFOScuQwI77L1sKeJFR/G
mEUnCINjbzZjSzQtf6fsJT7rA2bOHhv89mUunwtGX0WXP5CtzbAdBNIjTILipzC1ZOr/90iyUBPF
6x/xjM5wE9MQrqFMw6SHjrWFmjfEnx932/C6HE+uT2UAsKw4/vLr6MoxDuGHB5Sk2li1hnZLgdma
xDDEguJCOlGHueY7oNib8H1DnS60uvNb6Xd0dDIreuu9RCKfejgWFYELdY9ChEdvFqEbcz4prr1l
KAe4s7138MSi4L5fAT1oe5b1tl+uIA9O7+10bXep+gve3TPKweBVfIxayE2Kgsl1xvesddPe5h1r
+ZO+xAKyaPif6/xxnKPZf5DOniMGr6JHSD4gdbIK4xnO+jxKary7d2UFZUdmERnritPnQ+rtU9No
kITujjvK2cgtaMVi/1kthqluPyYIyKPUEd6VEzlYzPGJmkhB6OZOSvcXkJ5vpr6FyladUvlf1lPY
278bgKD/gEy07cs4lu7/807jHGdetJvjgz9lMdu7KfjxwC9alyZ/317wobm1N3IfZhKIXFbpM0gY
kp9R/R5gXkJCqjSGKNd/QGWI+4pucvjRUra0kH0cocqmNfI6b6Yw9ea9uVRJeamc10qpyZ4e++J8
52jpTVLsqnWaHYv6hywy//OTramrxo9r/Ur0RJ0RW7w5tyuiFhREiK0Krjpl2KN/lMjslsc5+iVK
B6zHnZqw5AAaAUBjl/cLZQ1poTg/JUjSWoTaROmE8oQzXTz0VXVu/PZVOdEe6kbncM7iid/5gDYP
9sOWRJN0q0MRkg212KwXjIpPsmBneDQcX8ny8AbsB4/CYp2CIguuqp5IpWZWLAXBWktwMaNpmIpE
L7x6iWpI0UXV+7LrW7q3QGOI+RaphTRbGTG7DRO4MfpxmpkZLEwcf5X6i/DO1gNx5KwQX6iPwAsN
VLXVDsGANpT7Y5WgSNOTx/oNVNDN8t5+91CHIP+UH6R9NR4fWhoV3gt4Tl97dDcvHx35exOe3fqU
2UWjNRqgH7s6FvsHZw7nvICDPFVjvVzk4oDgsiyKSX0kE1ZwARiD/tLqUJnr6Eo39gWbwnt6AMOi
xsDB3vf6MorljLhVRdjosz6BryTt+Sdxmvekxm78AjrIq4/zfAtZEARPJVQr1C21pmPetWpy8Yon
6n36nI2gE5uOk1drH38iP7lw6VC1pibv/O0535A1IVRAGXSIP3gvXmnCMsXSFa+JMdgQR76Z7kpG
No6ZWcG5O5zBM3QbqMOuKvcleZ67nxVVktZcEBp5JjLQ5VmJF+343x2OnhjVceRJ2sC0sIBOsYfN
ZZgaY9b4E8EanT3OEj6fcjpZBcZ+yxtL0VoSLvJq9ZqESE36PN1RmUr09C+KU0ABBx5Jx59yseDu
pWUcRB6n3wWkzvP7XqXzVTXhjCqetSlqXECVOrVQKp/q20KUz7JO1Tp3m8rGMVAS1Y8T2aJBh1ej
dC5onZRbyXgCHYruJ8pjwqC8rHsK2EtLub8wGm7K552yFjlkCDMLCxeGlMIYTsNdug9zufNdeweA
HOqu1K31MSKwXruyc4rIFGUR3tc36MvkUa6Uh+q7fSPiyTVeRROXB2r4yXF6cwpQnFAJUeo1dD1w
OVwSXshetzUgDaQKcK7lN4JOcG+zGytN91N1twuS5MFIqt8t4TW0yjQIvUJl62vZfhtOpBQBjtt9
FXnQAeY+3AsBId1rLWXGBTCyjoUg3QowVh44w6DWNbyPFAPA4pj7Zf/4TMQSm1/T1+6IRuKeN9nw
XZ+gWlnfDMsvvNEXo9G4nM3j3TA1PITHr8fjyfH2a/nO74mYpZXeaBQSqbHdIVPD3wydLYexj0bL
vVlmnlH46FaxAjoJrcnoCR8DGaaPh4REBhvBhUbbqZfJVrCl8kDkInLNJ3QVKf+GOfMvnXjKEVwJ
lIrhKKS1kHxYvzewyyFTan6QCW2v/GfyLSjr5MQOrYHydX0FliyJwEjVYzAu8Ik8dFd5SMmpDkWO
96OidRFt84ahqfqZGpG69Fo4NgYab1RIWFhf7/c4QVHoJ6QiunP3fAIucYW7LwNLUDANdwOncpIs
iSTubq/ef3ED3bkzkr9iz1Z7qUXyUo6CB525ED+K7+ThvpQZP1GlL547iGSCiauMWcM3fRSIrjKv
TEAmACl2tbX7zfA0PvOWYDuBwnxpCY65bCzq4gTw7TM1DTS1QCumSv7aGE+d7HOLuCDyxsxNnJ1k
l4MRx4kqQ7Um229UQdFQTafJXCyuwcjDwx7u3EhXagzb+ZfyOIh7eW5LHJiyzRGyWIS4Cb1OL1+V
yoR/ppK8ZEoEv2VdMpw/mkc8Hnxujv8ZM4VD4mo6s0D6KS03pwJPDmC3fN0B0ne3pKMTBmbjM40o
MNxPPq2S0dJwwka2+Xvy68/uzDXd0tMLRVApVu3gbayHZhMaD1iAaA9JEWeybsXLryggpCH8XD1N
Uqkk5n8/neAjjlwjbysGSoar1uofwaJjTRiLQP2wgjKWJC50XDKEoNxCbVoC5cAQYBjZhlxPfk7v
ysXFPVnHB78o/nmaWe2iZ8DVWDXdyN3HOia39YT246UYa3ccCI9gnZKq4T4/wqC7TeplRC2zk5Dc
Z1xblMezpLcr/9CYdCcv8OJjTBGXbw30zmSUOQ5wgOeuQDSr2x1aiiV+GvAUbW7YOynQDNvK2Q8T
QxMx6lkWz05xJSVaT0LV4CvPgdxeVIL3NRdLGrHFEi64ilEXFAIV8tpraHVTzrl0WdyPtXPxr038
Pd9LXxTiLPpv9iGlTlTZv80OhNHxG4NnPVH8p6Qj8Log68slZRM3R2h2z26NYVLfVvBy4Ic/mWKU
NyWl+MT/nA1OTwPoHNOW+ItQeHPGp9+i/1Qmxohb2iRm4KEWtTbKIDfZNSelNE1gbKl3Kh51bHHI
/HbSuGTLRy1NeASJfoeoIRMQ1XxQgKo6e+7m8BNd+9gD7PyFnSXXXSXtfpAndxQ3hNIu7xh2xuER
BaZUbddJAQlZ6OIIIlZOTnB7a87LTWntz7S+J2yokzRupPY6ghjCGatJqKSfx0aBwaVjpgdCs6RH
y7BE9Q9Y/otV1CJ6E7yqYTN86e07EQbrbtih4AEEmeFrWdNVTec0QH2PCP3YS719zhNw3OqLrlb2
xAmNbSWalSPhqUiVEkk4XFx7JRlE/FUlA6+oLsPRhbGLyQcG5b++MZ3SJf2Imgy8UVtWvL/OuDOv
STvsC/ro7BJenJsf+SeBQiK+NKECFmCEJxCEyb1AXj32BMHEYUNhwbv2BH4rA8KaVtcO563wkyuz
/7wpM4NjHinQLpsh0Gw5d5FfV8K9TQXmJEMxUiWP0m5pP1rkB9U71gAwnfdP3CopCT9Ee4Gkg7OQ
cPLxel7QGFPZ91elyznGYPBUJ7p+6m6If/fpBKMRv9vAl33HZex2MbEXg2t6k9ugemiqWR6x/7/U
QK7S6/wCeuqw0JFcB7MVcU7Gn8mjz9HNFvwxbbwtP4RxrTcpA/O623D3HNlPooU/mvSOTo1PkSma
e3jNE0kdaFdbyJVcPYpMu6G/rT0yRzk3SY3ey+uy/zv4LRbGEtNjWswDvle6fuwIw00AALCL74wh
K1FBF/ovW1Nww3PpSEpf19yJ7JiatnCtALhlWkOZDdtDqBj1ZzJAr4+A64KeyVl++izW2q1pPIR4
IUqCT4X7C8VtdG9OwNc4ON/6no/MLCRyKFX7hmqc/JcfOoYNUODuk9PiZP1SgKuN3w6iF3WCHYvy
51L3QwIIrrUEVL+8yUSBsa0FvhzTfKW8WqcDXm3h5PrkERT/owH0Psqj7SYu/S9ltyJ14Zuw0YzC
fCQ7ssSXTZYQSZhpg++vPTSADkhxD2cVNICvQwzJAM+t9fxiL8gAyya3kIAIQvdzbG9EjJcULPfi
Jn+0YoBPH+wG2MhlY7iRjNJr0MQoVgEnVhm1dFLJ0ibq2zjKhCVR5CI8uMMPSi34v0IaAQS6FmG/
ZNsnjw9VxnLQViw5lY//9yYlpLhqsh0Jp7nmknyOQGSV7g6UeG0TdUq6Fw2MSqUQ31uJN37jCd19
iMfE4Ul1RCUt1b7c3STI4O5NjqJmhVL1Qtvoeb7W68BXPS49gxXTDFS/llFyf9F0Ztx/MxyvD4H4
30L5kmOEOerU3xbUQzRAd33NgFFmBxxR7juKUwBpy0CQzTECTrcVa6dbmxDbVIX/XHq7RY7Ki9m7
Wd/CTkI6fPhlRjiaLMCfWp5mGtxf+Hg2lBc2TdLjzVmfVvbRra4WxfcXsm6u3OH62Xb86jv2Aujf
quRpJKnCyVwUeB4diWSt9WANwXACmU+UYfsVXccZAoVpUNlEYFR3SVTo2IcdXDt2tUVbao6ScmTc
U46JYMK8TPgncXYPAo1LlIFAx8845/VZAv5yWH0bUBnPGyRtDbU61ctxnY5Exj2mVs1RX6bFH/as
UCMRCKYSs3DandBTtJK7QKYMu398xVzLxacBWxr6KfpRZAYBZ6p2T3ixcZ0jkXpWQwKy3zrNcKyc
HB9SD/OCME4Q1w444kpMneu0LkKePlUyDcjUEtL7b8C6+w/PCUW5oyih4ZFZLEjH6h/8MfZBmUqz
HQlI628MHbmMx+bdOdrodzRthaVAndPibGXA8gU5rBzDWz5pA9zXTIX52ERm6oWBVQfjiG5zsvOb
u9CW7pY7kyOgqAQvEGj4ZhmX2IcFtfd9vBiHK4Jb8+8lbKmUHOEyHD8yR15jrdEh3AWYyUPIo/NF
Oz+7B945KU3wRvEuTWjk63Ve1tZihgWsnysUrkBvz4nLABd7ws0/5ylKEeavsOqC/iz9ai5YYOQ/
rWOzdL7q71CnEsTUgMjl4WQMMsmIQ574akSwieQOBxcjpBFt/fpZo05EzwKHjiqaU3bZQzZ04txG
XICEMSR/bfgrYoIWCMHES5VWkhGBbipptmjGlpIzU5fg00XkgjtzxZunt94BEgJT/9fzTikxUlxH
C4O+jY3U/aMY9nHxYF8vD+g5+J3ycBIsga5nItY+AElaoLb4pGMAIwVfv3vV/w9dc9W49K5kVZxw
T8wTTPr40/gWKqGQ8qGwh6UwQB6ByJAQ+Zr047b/gbSfFcnAMHHaml6f91YxTlzWWEVY9YXw8eMb
gsRIqlygwWcZ+MAtssIp5iJFEkLc1g9tNVRyUBCqb1Sav2GWyg9gyx6AJZ40843o8zsxlnjGrJGd
yw5WVNeE5CL1R09emeKnnHaky4C+Jclskwk6Rw4bdpVN69e5WrGUUU4uwadiNq9qClUG4AFH9/S2
xTaxcDIMCtsAl0Q4/9dfr1xAbe/nCr1M/FLeDF2N9p4zIsR9paKYVjQbEqIgWkDCxriBdpuBzC6n
nSPffpA5vxBxK2iUwbSqIPu3cu5TdqOWy8mDQglE4GNAZNqqj31tnl81RswNVBEzlCTvBOqqHg8v
vCCrFh3hE/c72UWz6TlMmj3DjwFOHvNBWDLv5BNQR5Z6f2nanW9+02dp3CEw9ppqNEvNyKU8fLAv
uKkjmYK+WosJSxjbS4XnpMVzb5CSR2uuCm/BbWyB1X+3obk3F0rFKrd/SZTycrfYdG+JgAEjArkM
DCb9qCIdMwkKTQFrCJIyR5txYfmVwsqhN61bDmvuIPA7tBkkxr1QVYDvpA2rrrDsB67s956VgUnI
QOTPtDjUqMTw2jeXd0ITZgAfDvVboaf88XorumAHOZ/nVXlizjQRHvqbyxIBsAJ2v39vPODgW1kH
gXGDbYmdZprAkkW525oAjoK7UFkWkK6pHLCB4oiU9V2G+TRZ6vnOsA+LmtOBkxCeeQFC4RSQ7GX1
pqL2q93/UtRTPFTJcZr4j2HXNnc4PE6Sst2CDE6MpKtiDAVPMB275GvbJUaFiBWD/m4MNYM4mq8f
iLVt0165HRUoH+weOT5CdWNR7gfu1AkNEkOh6H2nm3VkigTpPxh4obwj7JKEGiuytfOLVNKpPoWc
mZBtb23XGSvVSYenaNbkl5XxdF/z/SvrhD4GRH8Z20LtgTg2+f4tZ0drYOoUTgB7hEAV3GiOhGAo
BzONDIlDJbksK0gEvYKZSDOzdk99Lalshi0nMBRkuKbY0e2RwHMamTvpkyHSSNd9f6dkX/D3F0Zl
qhrsH82PWwLmZgEZ+DLJXD/7FU3y4oWmxMpNXxmAIRgRLfugcvdm/ZWOAfZMUYZIrWAnzUweHN/m
Hr/hk9oV3NsbKs9l9LyN89dy9Eswr9zLCv4gfoDks2CrxyFRlGDXp0ZRSvHBusV1F4OZEjEuh/35
jlOMggL0UvXK+bjXoeE0kf+yRqtEOPHKKKztd6ra/tAVq2XDyk0INlxOd3K3OIuXLUFLNFV+i6IK
J/kSZ5lCXgsB2C1CPfu9q9Is2BAuAFSDwiZuqMdwSKJA+d5Hz6FztHqrSxQOCnF1q2dRvNc6v6Oj
eEPNl2tD1pnJtq+aWoYdCZQ1rESg6mdszHj+Hjs/5cRf8cut//WFTdYY2xzl+s+7Isirljhcq0gV
FddkvDF8QCzlC0fct2kaY/7JjLUQ5VzfNOLCT4BGSma4RnaEhjahy2keTxsw3ULsvGsKUZzewTOq
oH8YHMQ6vaI9eDscykCs1HxoOdP70yM83FrTDZnOPH5k/sJI+MlIW6TQLnFSlkTmeeRyjHGvH9fy
otkpjklCV+eRSFqiQuKXqmrT13NBrEWiWLF5BpG7jUCfFlmbPvIDVjrk/ltbCh/XZBcDLcQP+JML
2uua6FjBqnF8D6sCECr2iOQYnoWx6rPrXTTNYy/YRnasRxtzivBHTa4NKmgcfkWP3Cpe+i2q5v7l
CuUGxsZEciD0vYWU85R1eTjmIzJ5azqBoxuju3PK5Tw5/iGuFpOAkHzoCw/RdQ8P2rSElJBt3Rky
WU2ykgQlcuWGpJpEA84K5fqPcBoOravHMW++JlaMiSeoo4bXLOofuztZEMN27LfENKOVADqIhdSf
HfdvRnjPATtYyYuCzlj8TZXrjrs6Jp68HukUKhnm2HAEBzkTziHkUVgkgIPwRrI0C6DgYTLf4GFM
jsFcT5KeqzchzXmwuTO5BphaTaln8rKgOCsGy4GtIdN2ZBpiRVJ7z9VH3NL1uISflg7JrP0fOmdN
tRDSrJIBp2KPt7YyckUm6ma0cYg3uoaf0LB6tltFwp6/WbdjFVG7pBtYDzHLrZR9paRIHucZTmrK
vpR8N7wFqp4jMcts+7Fw0r3GrzJX95ZC+sKcUG8HcZT5JesBBSNKsId+Vj1igWzZRkEG3Or6Z+qY
PvnN5giR2oUj6leKTIP7mxqNN9X6ttNXVh0GAvrPyS+Wlo/Mz9irNoEm1FrwWjbQfjZxhH0qtDZq
43Lp8l1jBRnbLGjtnJhOMao8wwYbY53gBF6EPNNlDku6Ko74fDo/p9ehlZ9Sh6ac7djQzHn36trz
6hlcAIufjhKjF5lFHXhNPK7LzvujlyOZR41Lna2SuAUlcVmSesVigmm0a1JpfGEPVi6Bb1LyzezS
dz2Q/oJAinll3iMZGAGX99DyIrn8BPAHg552DtgaaHgoK30w5D8Wwaurc/d9Dl6kdQt20dwrjCYo
I+j1ins+5jC2QaKpDJH9GCNWIkLTsnDPQ/f8aKrsjXxA7+EZu6Yeyd2oc6xFzU8Zy1QFOi9stNNe
+w/GSCl3zhNkyNppTziv50/keqDDDmgk6MrGSLiUP/svNykPPpTm7pp0ZX4J36j60k8jGLgIXz33
J2euS0kjtZT6PsOQKPDIZjs/RJcxIZHkZG/1kT2tLBIe+DYOAbi7/QajiRHIgweovzkRy5EpOqyS
wVHGDfgFqqA+uDXzYNL2PbmAliJnLy13McUea5bSF6drwy+87bGMwCKBYTUa7wFWRnGyqFuu35Bq
YDxHI/VXggSAwRHMzFbQayzkCj8cWGIER/a6D1CckWlB8iyzmZ0wD+19GHKJ9KAgFPP8fNM4xgRt
cTwYl8Q35b9oXL9ufrvwGUIJkyrlZ1R4MOwu/gPG8+HccieNYnsef0TOLQWIwC0bDxWXn2eFeDPI
ZIJMYORmZmTQxCiPB3UnpXSCN4uT/qjZIvZQpbAhHkLXuOmQOHAnsSIozJVkkbFWM/LR6mexNTLr
98I8Uf13GEEht7qfaTE2zffJSHnEcZkDZFu3NfsYU3LUaF2MUr6aiWxuxyHtnaAjIp/LQQL3eHgd
MmFjbx/nK0FUNc4lzQMs2v+JN7zXvfZGtF5wQA9SWy0El5eS0HP89U5qPiLLRcJazwpvuW99xgU2
oqAJF7gEbrQoekqe8Lax/A73mTAUQk8FmSXcPj/tNFSZOt/MVxooSXUua9cUHwXAZnYkt/0OyzRU
e9HHl1dSzzNJ//YDtDcJSZD/4FuJ9npy+ZUuZTBiaKJfCl6NkjQIspB+pb/cPJsaxxrxXx4MmgF2
HHwLAnAOUOFOFfIAs3dbvIblLwfIpG1j6W6pQsVSSSuBPw6jvdB/+OdeZRZiZMbSeXgiy/RpCP8c
1I77VQ8Ddkp8/M1WRwaqQb5lhCC1Nyzs6YOqOUaNaDGBMlQUSrR0SSmkUEZmSwI0y4qlS85wFo1m
L9Bk5OI93QfVj2StCewAac3vcVMlgXlE30UaE3Qwm3D+fZxiSjOP6hIKhxtPuNC7DSwfF/pL+ADT
A/CJtjAD67+vO9e9xdz3GYdKUSIqjmGrgBR5C+JkTyc2RrL6Wf5iW5mtjdY4FxSdXib/hkvD24FY
AkceuCuCOBQ0c5Lx2Kwb1cSe/XrahLB8rnV9QlSSvYv2g6QOwB3bjVzNPyEEc63jPpaCiPaJZqmR
CVhWPmsJbBVefgYixD80rkkE1d6uRVSpniASPKVr7gMqZywMJKIw3cPnivf1enBdJTrqH2xs8d4K
XG5QJIO8LPLC6NTGL8abgrDcDG56h4kKIX1jg0wXlZRmlT4RyagZRqj0wdwHUtzRXrtuaSAk4YAY
iKwTNqGCX8YB4z1YquH6F38SB+FYjAfAYyz9GirXJzht8D/MXqMZBzDadZ6DTssfoAjvdcj9Np/6
ZIU71Sif0WlQECLCUjPfEvPYQzVPdfjPRvu/5PeOcHV4yS2dHtzPp0yOWpBtmfGZGNTjYMIOo+gH
09xd59fDmjY7RYOqvz0HyL21ibBBSjjXzSwSnq6ycA/Y3qSMPZMeGHPs8DgAwOTJo7Bw2dYh0CpR
ftVGyElREpRnIRqlTw5oc2zaayMJM4BfokIPhac3lvAlEef4v4NBJlaQSUkjzxEC4QCyKxV04txk
1dGoVsg7fYI06SQxsX8nnB2ZNooyq7DiYvKqGnIByetDcAneNWYAdchnIp+sTHVE5PJ9KIebivew
MU8Ljr/Kpt7PqC1W8pNeRaHfnhz40aAdhY4lutEegeUOjiFDbm2hUHZJTDfJDnwKBoBQd8RKR3Mn
hK2ndaBuRbywlIZQHTEY8I+BF8rDmR8F38JaAc8ELtK6VTFkTe7tc/Cz0Brabd9fnPh/W8qGREQg
5Wc6jAAc+3W/sj99olRH3Rzuny4ZPb6nM41/LiU5LHLhHqmuCBkmWw9BPZvcUa3vh4GL6LvZVS3b
e7BpUvqn7BTAgu4RjC3sjRyJlQI4mwxqeKDdwWFfWa9yc5GxVNylyBMWNwzZKdkP3AaEGFUmPjr9
fWcSKR0+I+hi5OHWOquDkivMD7LOshSknmoUCP18q0ly8hG3tWvWb5KUkRRwoEojik4DsmrcRv+i
g8kpTEYRQ56OvBoyFiLaJfXY67cGy1hYWeci6EObSkSltdS+UrQwSALVZQqQ4dQH2hQq0AwtN2vl
qAX30TZEK74t/nIo58x/A4uSJZ4wwExF8232qehdGRxOQgQCcZpl7+WkkNqOVVgm7ETCpq64Klng
4chSlfxPg/TaZWaBkS8Xqryr0UMXcHdaEagryj1tKajz6L2Z3bBAJHILFStEnd7P46cen0DT6Mbm
A2zN//kI2dudOJMN4EnHDC2QiouohV6gVjRuFww0C2ct4WfKfZgqhQbsa/cZUzZSkse/VlVZssST
SerlgLIenY8pIoM15NETGLhkVck9xGMlqgbsvGVgQRqM1aFiPHqBk6Q7JhPWE2OCkA3amYVt0l5w
KI+ZJpOoNsIxGDZ1DISFUQb0M+fvlOEZIji7LFiAnGd0UceNDD9BanL06Iz/WIZjtrnPqYlESQV/
v6lM+KNFtGSX/IumOLiU4WRKSJn2/6iciMVKnDi7or4BOJodx8LR3/9Vwtx2GcpogLXza24WwiR1
vgNcdupOfljIdlOeu54sqRj/60b25cquAxOTf2eg/7wzMoxcsZkax2DmmIZAh9Eh4mBopBz+ibla
vMd3EmtthC7eRQMq7ICVavB6Usj56kD/h0KwwipQ5FQtFiaVgodD17VNrcsgf1ktNFT53vEqRAg9
L9y9yLHRRjAsT/xIyHhjLOSiMZfhTugPzUSxDB4MZ3PVFDIfkvF2cCUJ2tGl2ioivethaJoF+uY7
MbVl+cM11yGUiRsgjNyJyHRkHG1prlbz5N/ByBgHx4G5zbGvaYmNNt7U35+c4tsZw7T/3oNHlmhV
sOSThGKI8xcSIFe/W9LvYQcY7D11h2+k5qxMVHJZMIJJhHpUc9++tyqPL9Icz++jxO2umDVW7/Na
woCy+eChbNBJHe0SmL5ViS8ppiAzYe2a76m24MLoz3xMSLVcFIDAS2iAWl15HOMAIamHM1sZcO5t
Az8jgHe2O0tn/5/kt3QBnKDNYa0+Tkbn8ZTd8iedzEHOCiJ7BVPZ5EHD166wzc+Jxa8Y+Egd8gO7
jN8nR9EvkMonRDt+aS6N4HN6Jt2FCGKBRvqF2vSx+9VPei6mZYftIA355Lj3G8L7k+DYqLFNEagz
UX7q4h7SZZ4A1T8AUh2b7D7TV9oXdHi1VZfErugsS7/vxDgf2H+bajcVZvpVxis5TV1N+P0veyck
KHiRuANUQuNDHCtBM/neZijRyEIbScD5M4li38jy8NC7sdTh+hGDpT9bcAFgZtVZ60hKO0PhXE6f
SeUSr1OyuHKxTLiE9tz7BCSIE+LzsWOqMe6pu2gvtneLBIpmEryKcFqrVRf2WJL511M6vbbYSch7
FJau/FM9CjJb4qj/UHT99BaIXAAyfB8fAdOn8DBiXwq9XOXbiEbaR0/veD+OeW3Rdh2AGbCBWsJj
+lgTkLWcPYSEvN9iK1XbEJ6ZW20qF9xdAduAax1Rwc0KI+UiSrMFwXAxWNy1JQAM1Q6N+ApY2y0I
Jz2qnUXJx0QvXA/0eaKh6THsL7bjylVGc055m0GIM58LQ3GH05IXgEgtskcZKyKiwp6B/G0rQ22/
ZEUtrUhEZ8om8UNKNCZ38pF7v1XXWKbFm7FFRuOi9/qy5aJDOgptngXqdqCHFbGLhWrGDBu9rhgC
yEp+sHhb8FlGQCguCluTDUwA9L445ngeP27fpcK+tVzIlVy+WJTwrwp8j6gkBkPuaYwxn1Utl+My
ZBgiX+kIaC3CozcxtE43XT5zrZRM5q9fZb37J4PW8z1Lwok8JnhIFcb6sajjqTIIyjnNIygf88Qf
k5DCoISbzq/bfjqwiEOSHgRR+yS69LCDMY5CAydYx9XmIlPfxmpyNye0Px/A13CCuHcz83h6CVsw
7oOxA0u/IY4kt9JdIadsIIb+qvKIw98/zSJBuJ9gOo44DTrjNrIjgCBfkVZlk575JtEKKpnxhASu
lCcAJ0GXUfm7+m8Nwsk62AAA9IyhC1OJ3rT7jAjKxG2o893si99KnYqJLKgueGT1mAxIGpAW/zi3
g1ejAS6EQRcnwjZ2vOjqbznH9ktseEjJ7VgpvnpKSwoTTWYYQkfVWMqZxH6zkupt8P3Bt4huWEzX
DmLBRyaCH6C09AIfJtAs54TWfbyEsrBQs/DiHBpaZBx4SpCkII1akx/mhXmal6twnNaJyU1OTRrJ
40T8NEvcMyKQZJK5k6Eyk1IHeGTF/QndM1+GzPEz2+6u538u7j4D9gMxnQkFeSIdAVUeov8ssgrl
jp332JGUuI9oHNhgGzysvTqHP7ST2AZUkxgImDDXrRUpOqXFVNqO4OOVffsL2HJ1mrW3j3wpIk4e
7YSuLDsEgmFzOwo5f1EDJ/ICRQ5041iWCjoBFPs+1V1iiWhGMUDlpGMQFzfUbeABDsjtIOL/1eiL
8RJeH9b50RjYgHmTfBrKBaSM5iaUj4AhPuj4ywCAnJpY9CExWPotyb7xmnYyTr5RR0FDfPzd5/R9
m/UXPkmqde1kQYxlHWto0/Ts3hcDFtetWrx5Yi6760Px3CFPKLsaM1UshBtCj7kaxRmUBKpNdpjm
/B0c7xWggyQNTUjUgsOqqU4iEUonPFeP6JHtDs8A+rAJz0xlMM83XJf7M/g44Nzom+hA/SglXU4m
2BHIiufMlCeDj95SyJ8PRwufR39C1eiq8ESUK+qXoXCIiyOfxgDPa9vW2Or0FVvXa+sBlhSfK1CQ
x/orqWgYQwG46B0CEcwv5ojePsjbQpKyUWJ4VPRvp9f/VcFJyBtV16hHNr4TA+YQ8XJt/T2pnNX+
o96uxmbWkf+Dq9tF6WFNfxvUBmx2l1l6g96tKWKTpxOAWjnDqDIpO29PqIXvVZ4T4ymnYJ0cQZCG
u0Jgc2Jaae8gAQwDEvaXkrz8mXdAOCt/P+rEC+5/0Kvom2Fytxu5pDKWtKcYvEmFooPniwnMyi2N
UzmQWpRwetozhXRtQikV24SMREEMskr9+h6kkckNvxuS9hawve5TcjbRXvlEhaxEXqPS2lP+VgiM
TbMt7w7h9JQaNT1K9h7ojhv3GzMEMrXqjkw9poqALAUP3A6rbSzN70OYC0gLTBQO4omO4hJ3mOaH
bUY3Fw3eAm4cYCt4aIMct0K7Eb4hvbRnZeXvEOpVIGBjNmgXY8XuA2Y76BPgaKlBIFY89M0j+MsE
3HFLPqfeNXS2UR0hAMSm8crlfqToCwA72GZ/24tDzB4E18f7iwUU5mIwcrsX5Pa9XRBXTqKFfZrr
3dHagZU45aUdUUw9OEw7NmlnZQ2Q4VR2YFiEHY0lD3cFaZAGIOgR9jbhQ3nbl0nSOLamnUlZT/67
hwNT/1Ff7Le0AXeW2U+jcxWYx+uLBzDNmckqiexjD9THlrUF01h4XbG/EhVIDCl53NLpW2Ja75Zu
a7rVBZVsuycSYxQTjgBGteTNlnqxDTKc8rwJQBVH96MC62QYypFEmdFf99x0f8ljhrVFsMg+gf//
O8gyj5PBa2fRiOQN/N2gtq4GC8+a0LG2UDrocWNxiVp8Q2oH0fONZlR8CnffGzjCOE625DEgyDCA
O9YV9RGGkHU1Og65qXxLtxnCjBYes2BDL3Dxpa1D06WNcF9w9b87ecPEI0wmdilIFiN+uawYiFfX
d07GKGswYpat7fAPyFBJp51W80i2P59iOViFT23bW5tzrnokTj4/4zAxcmAygDuAmOMtZ8KPOPc4
QdFR3b78pZqPzI3cMYOPRAic/W6ssPM5URATVii/9nXwfzS7ra4LuAbrnUoY+1YhlnLMK6hH4LX2
a+w4OjDxZIP49SiF/1J0st5IaPbhVpqI+yFMOrKcN3V/rYHf8y/+t5m2XBrwdzfojsXMce6UhHEO
3Kbg2mW50hhn0R+fGy8bZV8KqJ2CAftFAlJKT7KRVgO8X2Cp7s5SYaGr94Q7yhs0PFAJaNobBl9i
vs3JIW7IqqLPieXVoN6fqxroJR12A+0ARyRyClSE3mxClJAj95dFiDBj0Wok7ETJB8Vi7BO1DdUS
NjTiSP5DaS5f8b76lblyMNaKHsUl/mr+L2syofp8Juzi4Vjyr4y4lha8Al8MpLxzLgNXwF7VIRfY
1oxjUThCL5cPJZJpH026I7BbTnlpPoJ1tKYOg2On5BCzyjlrUIMJ/xkrNvUFUzqo5H1Q5ZXaJgy+
TBOoIoLYmpVfKvFJkIR0BldpRsxbnhjYZQSeAYGafM/IyNXqK7orcHwMqGekecBLoeGrArYRwMQ6
z9ux8pZpMGpNpIY31zCVG35Xu21FtyEBuNDzYNiP/TzyUN7ysdKsS85n7tbhSJ/+6J9fR94eL0Q7
D4uBHcymoFkqKjCzceQ0oxVo7HLRk7M6X4ri3W/jugdJdoqKK1859KQnTx/h8zM2YJiIJNU1Dl6y
RBDltBDj+lPjB80yOu0jE1ac9OmROY10OymlFGS85GntOCZ71iZKaKPKCyyR82ACvpmmuUBU7iMV
/ndXB+2bQLWJDBNLIGa9Z1GQTbMcRr5mHrnK4wG3QQAopqdmcoZlEYd0Sz1kq/SoIQaN3zKEevtc
UsafKGQ+VJstzdwhNWEPNlXPbvlp1xbAYUQweqn88wTD7jCZEng5Szre4LDcFeqcq7/WUp8Fl5km
4j96CWCXOThkinwguOuscx2nQMGsrlRXB9CATeZ9vFJSBMo8l6RIV9szETeyMQ/3MJyHFlPqq3mL
HN/oO1eFBWBtLNJTIKeAgic5QHps5zYzpdSq6x3MR5d4VKKFHG58Ydj7mZ2SVrSZirJKb8hlxwGb
9/hhcqoLjAGdXEaw/du0E0hghhZ4AHkwtees5l5MqlzU6TQRv87Z9vZd8PIq/TjTbPJyuuQOGtrz
3Iqt3fuNyCrZeK+87f/S4UlT/zf3mmQDjw27/Bx9ozzku8P2oAUYtz/0E+k1NzHMcJBBcs1Hh8yr
nSWcowCZ5ivLll/DZj9RfjAb3a/5A1DBt+Pk8gCzvDOgxXypXxZtEm2ueA0616wSbLwKO78xzY+9
0+TH31rTRZAhqtphBCr6cH9DVNmPGpbbnRVnSe9RGnvmPd6mwyhEnq388bvjTykGpHAveSw/dZfw
Fl0/BBh6aEJlVpwB87v+u/ZM/HHCHxR04F7223b+gv8nmP7Gd28de3uk76KcstB/F1JtxgagF5JO
TXxf0YG9TNHvXbbjAmk2QXe5+7y3lVUp/VOsZEV30196zIyzyhVjg+nPruDkOEGobDLoy8xfEJnA
1MoBC8bv7BiSyvvigAI+YziUEHiRBjDfm62YINZvHI1UiaOZGb/5EZi+bM1UpZItTQq8NXHwCQOS
d6ZOF2Aq90X+5wdKhpUL3Dd7nSqjHkh3m37xwHBfOrFduJyeY4WmbKM3YKoZFwKG8u9bOMUMiRPM
SbcqRMA6k/xpkijqHe1AE2IepxMYcx/FRxC9h//7xWmHS09ggpA9YWE7aHdVVCrOmtykPtgrO1t8
/0oDjVdOAsfFUFMIdcGSjTvM9Io+7Kt8mBxbASE/QNfobLoWqkIT/o8l+Wct5+QdENPPItWxPNu3
Z6766fMeqdJcOKSXhEs9i0hKf2ocaS+cbZr05ZQiZtKjJxAFZL51I1v/loy6ugFjhcDZUEPfPVmS
bGEti+qBaiJR8IsKy4olPyVq6iZgp+gRUNtFawjfOKchMhwR2sW7Lh9W7w7zIqA/fcphmcnEX+cR
Ml67z42evSa/XL4YWgOgqsnCkxG+BkpWMqs/u1Pzt/D9f01fVhIHwwnI1f2aKQtrI8IFPnadW+yd
rz6I2fQ+REHNPMqvVEy81MSsdF8qRpRWmJGbR6qbkDR6EMOE4UVJsxh+8r0/QNTyeXKtln+374g4
xBP5lNn0uBbN178d5Pn8/BQU++MX3CbugMVZu1d1q+iLiHqBPgXUjRZRwOfQICAcSPGGP2+EJnIi
YNnHZTACcKQB5wga+wOalY9i+ZP+8ZFBCitqaQsqQzqWWkucCeZTDZDBg06C1GyKzERHv7L3qYkI
x4jRKPewPM45L1Cy1gv4KhlUsmJ1Wut0TS0U4YctvsKzTemNecfB2rzcptYSedutoGrP/ijK/jVB
EhrlT5QRecH8XyoKj2B0l3wgFT2jvlcrP4Cw6AzH0LJY4Q0UaHEqSnngquGKO0tl8ne3+ZOcT656
w+Omac+OTyzMAVdkiIjUVSnEnN08DaplsP7e0u+6wRGXik4ez90+jSg57ESnFMnOzqakQXmDzSwj
JIu05zxjohe2XOtRKYcbw/jbzyCDd7vuwWVWYegABcdqOuNQeNP6jBtXZDetCnPQ2rYsJUdSQrsN
DAckPQHTD7qDUQBy58sNZMiX06NfPjXlJvhUBmtd8fSiWCvWyVLgTMp5htnUIgOVBxnpZzsw0jwF
6VTPXeZqgTRy8HqfqSDWEeLXESrJvhrcXYS/7Xxc5jJ2TdcbZbkZziZFCdCn+Y5a1pOW+EV1+d0e
t8KZJdbfUASNZDp8X23zExwIg9a5py0XxlX4OQN1tz4DId0OhbCU1si2OUf0UBxkgWJc0SpV1pfQ
6xWSkEShGV8RiavIvPDTUmhlxrLLgmDpck3U/9ycOnpJltyiiOnCYyzFES/QbQtoCQyWU//+k9fm
I/MhZSDObZvmc17DBDAiues4HLDE4TpfXn5B29/SqWTnfU90Wq767am5igN9cw8j9QPFnR0uVjj4
B2lLwh2bracRkRc7o2AUY6m80Ru4EGKw+EozOBa+zmqmXT8Y52Kf5+yxJncucRoOQALijTHi9sGL
9AkeiXV2TyjKKshw/X/iumOg9bbXDHZv2NmdUUKdjTs0Pn8K5TH2NgljImSLwxJdi+Uo85HqUeZI
jwOJ9OvFf0NSsdeJgv1IuyRvAUI1TJTrt9FRzSYmGSfFSNW38CV0CAeEwO4vCAbAoXbq+uul7JgI
+OVkHFYU/M6XZkGF6BaxKmyUb0h6Bc1/0ZKcPD6iJuaz/+YPMNMn5GHtEWyWg706qirSdwY5KP+E
15d8GYMRUqGveO05YfWaOLt14aa9oas8g+sKbyEbcPjLgfustdndvTZ170VQI9GLb3H4axS2tKO/
DKf41tiGQH0FBQ2sjEIfnC6bGSxRI++hfMTm00Xx6mztbUIlQFZdmDeMP3RWDKygUqYlte81pyAb
L6XVaSF65GfvjArsajW+/ScP5RwFHBdzGlHrGeBKzPizztN7QxhTrzcdwmVOlYTXkaQdJpNvQFbx
tYwWv+kMq5obROIbc0mIrecttSJdBi/LyD7DQ6WI0KHkENrLG2c0DWOnssc6InCTYtcJzk7MYByH
YMOfFsMl8BlM8iD7TCbxUaULOixYOIyADlhdJ7iBnTMU5KOmfNbcfRmbKW7BYrEl1lyUQW1s+2hv
mVuLwyY5qtOxjF612p2egVBr4CQiqD3TKY9xqcemxsF8MWNnDSIv0p66Wph1ctGGCVdjemBqdOmv
V8AqBBp9LZT6OqYkE6CQ/H5d1hgnGPQg1Wopov+kKs2F+vFtup3ZHx+HXtT1XcO8S3Jvwr55z02p
xKzDJ2cYAVswsZ0rMJP46DmJoeCujM0TjxK8VyQLmNsMM5OLTlVSWIQLPcPdppX+zNqpxplIRm4k
+Aqb2VzESWGBIkp9PE8/0JnHF2EtLdw6qKNyTK++OSO4ifWNtC/VdKebkDFFSbZ1LCQNVdsc/c9F
ep6fc4vgb2akrKXPxwmdIhNcskRrNhRhcqRxACtJzkDGRuAyzcA0mELM9xRN2yWlV2/E7TfCw8Pa
6SDREfRBlN5e3xwnXIs+7BNiGjjH6Sp9hmOUykOhQaIfot7zXJopdnG6djuOZ1ccLiJ7D3s4vlWj
gdW43SoMoxxvC1kXy9LxKBgBwuIjzs2qWxvwnJ3No/AVTIDgvib8kEPx78nJbKl3wfP2br1AnUUg
whDofectTRMOmUMtixTMc4PGkueo0x7JHSP595NXxC/5N6Bl1igpJUhD5jiUk/UPICHUO1ON8Ve0
c+AJvqnNDzdjwoW7dzrOMueEx9hWjxvJxfcMmkWkzhJlswf+qBgUrJaFfm2XHkNJQYbhZBQH3gZb
TKu66mh+CQgRBpR7pXpCcfc7XH72dvsfHx2dDqf1x90TJ5Ungh2HjbWFeoGQXMg6/eezUDI0l02E
1CWsIhsZRsWFSf69Z9KK0MWp8ugnvYuqiV4gFNSCeLpygvKvjmk9dph9adMaiX/MXcUyZjkgJHwU
oCj66OLws9gyZSrJOhN6+tvQwNC/KCIB7nF9T8R9WI7UleSfy4fVgpvStNpmAs62TW0e9uL4Dz51
cY+3WtRss+LsbzPQBJBEa7oCtNN14s9Cl6nYQa5xtdQGDsV1tMXT0aeHemQMl24KanaSq/xQk1fR
E+dyKfquW49kEqUPHL9jSpBwT15vJCkyM6SC1TfojJMA9WV9BcVZEBoZ04BIM9gzCwbzclW9RhMk
a9vqJGnwhzp5JBrqg1CMgM2tvOkHfEWkLZ/2L72eyn36f6X7I7DPt+opM8bfmJbBW27zJCyu0o7P
7Fd5D9sH7m7SRxxVc09ICMQx1nAktlyWLjEXfHBWDL6YEBbN6sMs39/nt6TmDKETbnWH2P9CLOGi
x+/WWenoUB9SXx6RLI7NlmHlFAAZMfn7guRp5gRROA0ty8ADZMRsz7uFyjf/YWuECXy4P0jBTXFL
9briRSkN+WzHBYdLvdD/2aJ+PlqfIczdWKz7YQTW56Yxc+5R1uohyMQRSx9djrRgE28B7PuRLcpf
r2fCFT1z7VgJXTHGfpYA4bn8qI/EjwwN1SuC/3JTzuLyuR+PhVOdFRxMEUwpOgt1P2GdY+BtNHNb
R6gai3G09WVaIAVK+QlW3xKiblsFCrEutroo0i0TQ/5E1fxjP5uSpERbv3bZLt2Hd76X8pfAzH5I
z27UO94wtQ+y0dXSrt1LHLgBs0Pj2e766Qqy9U6jchUF6E69r97NA3EIJW2HS2Gwwyphp9FxrJnx
3Jq8+GLMK5qu2iohDRiFgcUd+VAPXl9GDXIEfmg8RO7ocgiMOH5v6+FheDOX1uAm5BIDw9sattLw
FHiebmOQXuxlFviCqLYfU6FMIrMpJwmJ6JgL5FO6+f7QQIW8vzxzqtM+1aaX7k/hHW0pLc+YToAZ
MHbobtIpvQeMOy8cN4X0WoRHgFSOKB8jmJ6bxWqQA8AKxACO0g5fG48z+c+PLLWKfDWTZQj17aoC
l/t0lN+POusqe+SxW8T1LedI3h58guVaHT1q8PM9h8VQk/Au2lBYlUvIQIo36d2B8CMe/VXB12FP
GjUZRGbk+OcAkZW18/FviJMr3p1Uy7MKNIePqGZKZc10XXzpRCWeLHRQAzQfDWxxAZ9u9M1KT46B
SGO+tL7j/Oun6bcXRo3+0Rf9MS2MOqfO+6jMtTT8sm1LFp7Wd4YT/KIkQfmKxjke8wPyOOqnmLuu
+1rtpUc1eDbQhgGZ7rhDT+H7modiP9fvb4a9oejiQVtuLWkgSz1unh5IkL9UQmgkYYKhYU7SUsei
jtTfeJML1w97lWdz0JwLT8K0hggzdhbLdgymWF9C49kIuJ/LmYJE2IsUTDsIJjH43mrHs9ipPQ6+
HCaIEJtsHdGjFyTYWUItg1BoWfxDmxEyjvpasXPDvHLNgdVK5FouQk7i32+wTUFNKEG4XAlK58zs
Z3baEy6HCdjTzChaJWns6FKmyRtqanC/QuNpz630pOyGHNyq1DpB8BaXcyXzyNhnoDjw0iBMnqt1
5IRumHdg2d1A9cWv2Eqg8HjT4U4VjQx8pnyG8En489PzR19arxy7mPb4Mz+xTqE+XMdz46c3xiIg
mdkBxiJnoX/pfVuz0OFbnmqqNoIlXAu5aQxNFzafERCQTDHXv3r/pOhy1fndbAslsLlN9ZmtBkKI
wyPvpSpWClnGQgtSY4r2jjjo64x7j9HAyl1DRgXjqQ9jNsRRM3YBzq/1DzIxslY91YOx3wWcS6WW
PxM18gFyhYgzzxhmCxKoFnE0r3s0TaVEldHFpVcStSSroBVCvhcpbTUXX4n1ZjxWX4dYzmXgHub6
m8jJm4/+XUbD5dVsYG3+EPc0aZ2grddv5IN1rVKOMvDGUq41w+kIhrCC7QUMx1q2pCuCn/u7f9bC
cMPZYQFxF9zifvXVkDQ680EOMlrEqa5LBKhUcUzlvfHFtCQyprEUK9bHdGiTpPj5opMKpXp/wyUE
eJnkE9Exjzl8POFKqjzU8nBFsyfTuoiSp6VZlamsOansu4jZobaRwxW9XYKdck2PbAlu+/bw0fwS
mItjR+DTU5eAirw5e7hfdQ/KBSBJZ3UJ4bBqEp2T6RBoSJ2C0OPGsmRhbCE2mdEPOwvbRlT9zb2B
19c4XgiopTkHzmwNV4DNFAgV3n++5LuLDviM5fmM0N+P3d2kg0NNlCMIKY29k+Evybo0garPC4/Y
2Ue8LdBuGDhLSwyBDB6bLdM0/UrOtmPrDEvIPl89GhgJmQEBoHxPGKVjmBsQgD0288Ki2xDd/zGp
kVezksRAvmm8L/loFezum0l1RkkB4Vb7c++QAnCZv5wNYm762XUKCR1jO+MZTd4e6cXhMfgvSdiS
BspaaqJD4CLHb7tAORKhhKrEZ0WSAdKjETpSWZWrCvNBuNoUQojD/eZia+UztTWoKyIuPWTAPBSu
Lo53JcF6cdFytB90t+Z7BXxYEBhktcLPap11NZko2dt5eJIb0zzcbeRI24KslxT7alkuhFF4pEp/
OO7yblqstJHGFXa1Kyso1bkc5uK4ulozi+cIpzLqZmvbTv1Fm8tOEsO3at7n1XZHWmzw2sIFmwgU
WdCdPSKBhVhvPw39NcnDTlwOcXQoqusWd2pxEfdlM7bIL9Ml7eERZGivAlts8PvCEeksbXoCOWlu
/2j9yNIe/AXWUebVaV+r5Ma3ajl9PYJ+Mdr8OqkGH29bBMVG4w2f0dAK8bYpW0NkWkcSHvKXiX9Y
sTbMp92KqdsESc7NsQKPMFd+u9088Dd8kF4TbdCFliP556u+miDTUgbgNg9p7Ybj4K1fa9TbWQnb
Xu0E8JoZ7Nm3pIUQbGW3Q4UoJxom1QOyiVZp70J9xXTtnVSg62PIx4anvSen7VPuj5OO6X4PTpt5
/kUgWJjiFm0gpNtdBj4f2LGQpkQ+M7A/tgc/dnocru0gz7Z2Ao6x4PH1y5xZju8DR73LobTcvjWl
xo0lIvwjxdPFKN6GqY+5uT+trNn9UFuP9RtK6CIDQunIQVkOIB+PWzGpQMGOK9yeIxZI2tnZBtm1
qBs1OGtdA6LvH86QdBXPVobwJul0tnZ5hSiDJwwZxlMJW3450j3x69zSCYMvyufXfRG3tt6uSlRh
GLKC+ChrIeHJUcCiVrLrRX6956OvleqxVgpbuthGmRnQfKR5NH9cpxXXIfCtpSx8kaPJHRCE/jo8
0qTDSr0e8Qk/VlrD5aOn/Wodes2/CDXhubxIrotwiuvK88lvFDYMgmxYQYBH5kNucBQId/lsn09U
PgtSnb1nMjYIgrbFIRl3Urqmf6AtSoSOCaM7OyYByJwc9+NWZpgCEiFW1RtHYaEr55TXx9UaXHi5
IAuuz0iD7c+rlerH2V281AJYVz6GSq3tjnasAEJjDG4b3gZqIAamEe4gojmiBYnj1q4hnc0GEkFS
Wu8kbLAEGC4HnCCowWi5yYeZgEDgQMP0VRWhAY6zZopSU3n11GzbpEKojYlrQTaTfqY77iMhN3nO
B42y7IbS5+eU/9l23cX8+45kwcyKIeyU0kZpEiwskMMXUGtuYCWa7tEIe49GP1ONdRcP+6dNq3s+
B/J8rwlqU/anShHgoVVxR4gdkQL4MG6cl8+H98UqYc3Mywh95829gvwoOPFDbg0JfMoPFyDFdBp4
1KyRBk9lSSGw/dgvJR5u88MzJnKf+kowCxAHNAN/bq7qSH2zFCmC+uinPXCJ6gblpzFh01uR0W5u
0ojOPRzE/5MNuB/4MUz2phrB67V92ik1Rrq/YyGA/t9pdULVvOyUb9S+claBK1qmgmkKVKUomhV8
GOVvs1ttOHfr4QxI2YKxZgthconQF+YI3x8pn5pSq2ESPvACL5qR6YRvYLxQfzvu07wrIIHEpxai
Icj6/GQKe5YopklhOgj75npZwtxIIhem3oggBXIX3H+a99PYfESctqQ1EKEnOW9yeE2uwzfS+iX3
aaHj3pi8aX8hwC5noLhKlPDV81shJAR6gyzO24T1c98ZTV+Ys2OM/NZm6VLSeRh71eJfHek74NA/
HfaiqSf4Gg2cyvQIAQEnPgcO1N/T3wytzdl6IQNsUOSru6BwojKTbOwcnT7UxMwsDlKqEqWGA9QD
rQxrWRqwHxlmY2qoj6uONDgsANzjHMSvQivjUt3RKp3/L4iDWWZUG0by/me9SP1mR0oW2dncwbSn
tMeCKU7uycF+qsMNXlZ82dvrJgV8fJUMVsKCZq0jnm74iT2WyMcxLMk+zDcjQ4z4gzjPot7aPfSP
fv4OgCBORSdiirhuPLEIAQ3afSBpK+dHOrj+r8V1Qz9k4QoH0+qm0tV24MxK0TT01+Df7psZmlTz
gz5rCwJPhkI98GqUXdO+xEC/NX4LVAzF5swwP9+j/tVH7SIBlH1UVfsKLE+h7dFAqLxno6nCpL5J
XMEUT6c+APwyRiXaHt0ZfBH8ub8VWp3UU1+yPIgPI7svDgd9eTTdF/vugt8t6rVBYHcl/lKbHmOs
nfWijv+frRfKWr4XjQng+vr+tqOB7/UjJFlZofu2sDihi7TrrZXM1mVer5SYsJXVg0eU1xmY71/C
Ad1X9YAcomVg4GehFbxBiMCFgPmq+1WEi6Jb1Wqj/5mx0wdpbpLgk/GqpmquBUsX3YWBIuOEsMgB
cb6+7WECL8RlQOLNFyRCrq9HcuT490z9dIqy8S8G5z3zkMRBWAp6K+hXzuWETvAzE33sNCrcm8/z
a0jzNmgSFZ6lO5YU+l0R6H46Hw37hGBxGHdV96/4JYnMyRpM2a4zqc0Zes3L4EXEJRCFdpK90lAZ
/XHBWlyd97/zOShGBIFSgWe8Lj/4Mw4F8NE/lnmjoQTZFmtiyp1b7WXyECGRfJn56Y77D3WDk4W+
psf6z3CJcQbTx1JIsgncFssUMQO0ptvyvWkkAWtdoccRCqGpXscIIE4nQgzCWqQ4A92BxIjvyqHI
6ltbcvGOutMmZCGRD9tm1EEf9kZpea7//IAzywzIFiMAEJ8NNbhlB5OOGOUyEaYh6sThOqo9hPnR
nEuNhGI/XTuCYuzD6QY20uukiLmLx3XcONosrGExPejY3OdSgh8F/8Yw0Pwwwgj3Bkh790Sj3Wcw
bWYQM0jgHT5XPC7tWkaiVuI3HR9aQyLTczVvkLd1sO1bxPE6sIkt20/T7l/ZdpiOeMuprrJT+2R4
1tAxyI3XQb820iuMreCBD6AYjU36p0cHR8A/ZXW1dTY0NZ+8bwZzJb/am/g+msgJ7jph54MwYbzq
Z4X7RTPSC0injVARUa95oADiNpOUwf6iEGcQRl3YBbNPLj8wX2dyxQAX1h0OGvlzdoY5b4eAeefk
SbADf/2PqngRT2lCdlanuklGig0/zTmrdprzs9OY6puTWGa6Mislj3QLHRntT/cPREEZIr4zonH0
EOgRQO4RWvDdGF/1prZmijJk+l7h2ybB7WLzAs0/VwiFuVow4MYw1DWiyDvKbiNnsYgzLeB8sriQ
if2U8z9MiT1DevxVb+/JF2OR+eG7bpJXNahg2BL6DbL++cOnesTvIG+tD4XvRSiP4V00C6aLDPEu
R9ya1RCRCxc55xvpqgPmVN+MgAx2hXYSr/h9zarUKuD+9fS0ig0CqjbIVKuLhWttNZTbBaqi7Du6
bKVHvmX2dKxCFmkAt0X4UI/FuprhJtgce2KRwiiQkjExSJyUcM46bdwVU8jBtk9/WrjgO6Abc+WH
Omvd41TZ4OCXC9Ct8M3VQ/1FEMcpZDBGJnZ/+2pCaK0pi2+UJOvGI2pLTglIl3hCyD/U/f9uJsPx
iWIzxPHAoH5X1It6HR0rBNEp/7TH0ys7aH3cmArojxqpPZ1hACV9qx12neVsYzt3PunmgJunF+lU
ktAk6IzURAyNgA8OMBdB6E1ZedXAgObvVNJrJ+7X0io/Mx6Fw270LmLl+Vq8U3xF7YIJT6QCS3E9
dVp4g6/29EUxEzdMBm7sFmkY22JoDDnT0Z8Dj6Th6VlTiv/CcEdO268a2t0j22C9lWF7ekwUCoM+
zPplXuJACo95gDwx1bqgFNbdr/i8FP0HkDmIHipBcWcXscu3bEVZwdaj9lwCmI4C7ohZ22n8pW5f
sRif9p4R50X2xH/Gx9YQByPqucoXkycCxxY8Z0y7d5tCgItrBKNErDzh8TFMB7lc4c9+DlZTUpAc
i80ND3NQoNYx+HSLsbYE3nNIJtR9Y6BwhZipmQARRJoHYavWHoiOcnPGtcc1eMDyp6g3XGcbAhCv
VKiqhXNhCj0W2SMUBQtyjOayM5xMhWVcHrTemY24HkjQ1PIBKZ5+AEyzvtU2ueaZVXHkvvh4z1KM
/q83nXqdSYH3LBzQOGUW0fzrjVWJo9f7RL3u6fFuU2C/VfztCYIzDSLb06tb+S3j1vfmghCWdxVP
2bd5M4envN6E3Tl1ijZ/2Qbkg9DzpBgkstWlAAVE3tpQFjKaTQ1b68eHZuyRmpPNR4uhcoM2xI3Q
0gOBG4N8YJVQhX1QJ1zUdgwfUZXu9nAb9ycEcjkA73DLsc7Rr7ovl7js3SWxeoueHZD/Yh/OPir6
g2VyFmUUV9UlE9Qt+cf+/vwmn3IovPtmHriqaRCz3O8Md2q0xUhlSet1ckbOFFyex7+pISF9XjPc
h8yyhQo9O2vXG6Ai7+Ij7y2SC/yzuXaFwgHMtyF68S6w0tc/xjcDIfToAqtR1bOHLNHxYC7FvzjT
LDJgVNSPoKTXK00eT2mEo2CKlkSZ8GyvSC4R9BlJNGHlToDOHq5IFYKq/3bav/c3ITT4INDHtE5N
fXmYm41Df9CWACTpYkYI0AFML5EIHzQvf0poDnaZgsJaeFKCOGTPpu0QJP/sjsrACjiRfBo31sr3
1SOsmyDvGcNmus+DuBXK7i10we8NCzxwebML0Spq0KCdfV9D/46ox6sZJPVqh3OWh3edau3RzsE9
ZwYZZdvi8j90rnpXr3Xk5FSymZCm57ev0bVsxZsQ/xzaLlDa/wWEFxIfQJkvDEPgblFI6uLyqv6u
4pa0zJ9oyp4QZT6UGK5uU/Idd3KCVybAEhZPFIQPmCYmXyrQW7fIFiL9izaeSB8XF2H0i/xkpdYj
ZI5M8bUXHabV9ZXuC8+3UhW1j46xmv2a2PysZGdCFNydt/ND92koxP755FwdiVHKt2aZYF0hM6Tt
yoGu4zxdKcwvd8JxgyLDTBFn5pR/Bs7kCjgyHRpskr/00koLxNE6wmM3IlDQsSAHiC9oqrmhbLMv
HA3zMJxOOXGtqIULSw7zfIWQrChSSYMfVqLlcmQlphb1fTQGukbKDp7TdmgH4epqzq1GS1Ww95ij
6WA8j2u+z/nHYWPpA81fgXy2e1qgzxFFd+YDiqEIlHj6AOK317W5zY4cyWULrW7Vupwj21aqMNnm
lEEWKr8uzX8t8vRZTABdMIf9/qlovOmroeeuZF7RD3XzI0fRzQ2N+fOSsrBFraMW78iAEsAyo74/
lkDRl7ajw/3dhVGNAfB9/UcE1EXRLUaf+aThBGB7FPKd3j21a6zDAbGjMSB3MLeb/VxTUi6Pyhck
lps0SxutmdrCLae8aKQuyJatYmA7m+MHnBzDMnGoDXKSBMUKBDHhFerOCDqL6sL4KNHRQTJ2ezC8
VGtlP9qKFJHUzADDCbTq5OKeMXScUE4tcwNMd7cyYyM9qdE2cyTM27clEhdfQT1RfVJki7Ov/VPA
hcN3NKVIIm/O1Zqlb07YiaA4ZAnp6B0ZkCTrgcQYvcwJtY0lKRw63VYGoC/i+Jf3GyUbnDYDidZO
50tddl/Vet4oP/7Gu0PH/cJaDjKhx085rYJHGWOKxp8ostBerdDF8uEoH1GCuxDuKsW8j7xlz8eE
RTZgVRI/0JX+VK/aM15gXlvygimBHjyWVjiOcov905Ss1uHJiBeJPpqUTolRNP6eC4TJeHJlkama
e//RGO6v73aA5ZS7R2FT5XgOPs5UI9ub58bM30UZplR7rDSxIYLxa3ngN0JDLX1WkJKUwzlE6N/s
gfpClF8cBeGxwIuouNRPEBQP8F+M0Y85y1WHhbGG+9ciYdRCsGJyQGgNHqz+BrQDPw2oPlXZmbo4
pGPK6P9Vmr9o1xtZ/7WRrpbqrjSLJV9szVL/nHpt12QtTTl/ApQ+0xtGyYbXOiEhIfQGTpWBRQBs
OpgtlnUqYtrPu7DhGhBkw+gxS76VfeblPWUswSd+TuIXs4W8aWmA9oAPOjwLM6DD+KeSzHUtd4fT
vg4jy6rw4gfcqvR4eHiUcjya61yJ/9+eyWCOh2ACRT9xcBpQupdcBKK4gmdTjAJK3hMf2Y1YRPMn
BdKGA8J49A5OJLvP87EIKdHEPygMO7dzQArA78D3aOWcT5n1uQ7DgENMyoRoNNxTicUsD49mYHKS
xgWSNwooBu+T97DstRDhXAkxt9slne2FCyNvyzBvSPYmEkGoGer5nn1Jj3OoaEVaBrtP4HyAlvGS
Rd0fow6KHpADd5CHTK462y77Mb5xptC1o3ti3MtnACiFjNRgCUDqRgkVwCx7bnti34AaPjlyXVSq
JflRVx9hlkYirDsIdOj4f5biJgH1gz5AmG4gEzACse2e2TbBinLYERV3z9PPpojUJ9JZDPJ31xUO
HfL6hx8q+fF50LIa7kiyKAJPzXQFHe2xzCBPV7A1YLNed/FZrJa5QaQW2aDUUlx3TcGG6eizk+Mh
oIjRW+X5Pq7/FVR1dOByylm2k9gpk9s8SC+8S4QxotHXFzPr8dHHEaHLmsL3wsgKc8JP5DJuFCxM
TMqHSJxu0jZ6a0b+D2zIEumcRYFOVN+1biheyCYiUjn3odcmCpO/KQpnerSbCnadLz3K3i9W7hpe
8PbSfB3cMeelUrTMGzHWklIt0XBJjgjmvHfxd2ajyA5yi40Rimd/0kGGd6TjOhKb7yM4NBBb/7C5
/qnhH20U9tOZwmW5CAG7AStIGTm6LExi2u5EWoLOfyIIQ970trWopDNgXrmYgcjYwKAgrqBN4o3S
d+KwTogkdeE/Yeup/3h2b3EP0M4c9FKBn3nnD2HMPlyYgWmY14Pp1O0pIffgj2W+PqIg29+zfGJr
fM3KIf5xZKIdWtdjTbtOMAnIo/21DFkOY5/wHk62npuTO/X4qTsb9/y+3Ic8uHY1wrgn7E221FlQ
PivfkGYvO9yWrtHprHxIMjJEROnvmQjkXgRH3ILsEzmbM0Mt2yN2/QgCd2xHkJ49eZiAYfh41n5b
f/OSxzRfPu5khFzMrQi1gaGidinyJfKYPhCsXIPbqO8seRXFgq+BxPyF3rJDzr/hIQeFcIpy8CAi
1xKzht/A8K9ADmADx6epm9yNbrpUh6wc6M1OhMhmBihQzO0L3ElQxngysQ1suI/Y7qpxSQmR1Hoj
7ye5GWodn8wsyMGrg4HbFiHf2nZYQZSZFObfPilW+QbUA9nOUFxZWEXyGak952p6/AWayG3pPPAU
OX5/4KOItUaKMlC0YlVM9MgAjOno7fRDoEnfrHp1G+CDRRbKtj/14dZarbgLtItthM49Z1jkofKx
dMqN9P1tHf7LtOOneQjp4+/F6sntBjurdUMm6oqsvmlkzbH3JWZhWmrHn/2u1LlRznIcC53It+iC
jOEOsP/P0+mR0hfZB9j4w0jbKJ7Si+bhy5ZBprAJAEaw21YZ7BlsVziLw4oKqHx2hVz1Y/Qf6Tmd
OtLYmryXLKIDyAbD9Pa62vXWOVbHne9h7iiBbs/QJXVH4S7G6/qM2l0UQ5C+t7KsUMFpClK2cRRf
GAfEj0z27iZUSs3X0+zeL9jZkmKi/tSxx3psNc5zuMuovzHUJmzlpa4psUvrjTXs/P+RjMwRspcm
W2b+VDTPf9Bdqj5p4wg8HIpoj/cBedWudJ1J3Wcf0pPIe0e4/oBjgJiCGO1/QhHua0AFDAab2G5k
34Ihgr8pmd0uYYdaWn5cNoVcbhrf6PjritQxnDUE/B7cBFHOxbWynHqwdBIrcskhu9rWMnm2RI/k
l9WMYSWwhYO1oN3o0kDoPk79rZqlxZNSyLgHQmzRClIlAiWqzsrnfZo/gZEn8pdp5ONxjoR79LyM
dLFM3Dl+JOCmUBZiynuh6Xk9eCjuXm6WRvJIJ7gXtHWG5ouoXwzYXvY2j1oaxJH5TSx7Slqcq1BO
HQiWo4BuyGv1uI+qjJr1jlHkN5N6e4NjTzmhr51mdfTmhNjxoRVzv5BuvUxba5wgeQXWzyuo7I4d
pEwJ3chHYGcHqdim6O0PJ12KAWt4fFMcgeQ2J0M+edR/LAs+UTvYoATi/Rn86exMeqPVPlVbmxN1
Q4lSctcnKUbm3DmZzPKRf9sEyzSr2f4qlQ/qkdOTwdZgmdOfJAiJDIKMiEZUnHCLvzc2tAxcVcHY
36i5jS0IYKgq27qDyyrCM6DZsYRtscMYUzmQCtrjMxIs3vlzoEgaiN7rFRMnjJj33z7RnUXK6YEa
ZaSlJP1ycHaW3Mo/cWCi3mGVAv92imMc0rAVKYtFBTmPNyXUABO7zwkFiUoLu3p8yRVwtLiYOmWP
gmSMEJlOes6J3Yk2RPue4Pk9zxPdhYvplw7yKWO9bNHxvq24QLqTmRAVK2V0ibAHkLNT6jJqH1fN
DKX0cFV/eKE2vhFXw+wZNQVd4/vKGxgo+EtV61jxWu8XvNnrwNAce3eplCrjQne1pJwVziJLlWVy
vY4zWZ2M33FyUwfvYIq3wRCFoG5URDenIN+pbtIPJeAGyoDYFZ9NVYnspX6kTU6fHG7k6KSTf1Qy
4VLtnC4KoBUuK5vqbL5q154FQ7ZHEautmTaZPptVjL4Y1yUChMQmZudRAtwvGe8BnJ6BiLhAl/MD
XnJCTSpvHR75UFezHpMgm2EElsPUQCvwH0/dineWNC2K5YQ0faHHG2GKFZ5uV8FnAEJMDqBPXBQz
4GAhhWlF4ZPv0xkwtbE8K303OPiH0yEdGyUrWYEcW8x4aG/SMIJQnz8osXM/5F1vc8yxfOhd4STW
WGEp1Eys6gadxE6hCW2++jUwOWVRcTdB7XzNrRyPbxHRF0Hgl8PG/EXnPSPF4PeHfTVKJKZjZMnF
FSb5f07uJEAq0ZT4fw5Grrr9L79pzpYWd1rdNSJI8pW2y+Efr5uCzrS5nbZOdnxkp0oYHLjoPl+3
V3ubUJnqH5HMuNuIZrboJMtafZxD68M1AR4bNvIypsegIlPiGEpscEFDE0nakXeSV0nYakCoK0V5
c+ue9H61mmj1rBK3Xpb9OPvL/wSb4M/F1xjpJpgJ1b9OQbprGVt/R/n8s9zpf+A85w/C0NzOQ+i6
hxzk5nw/qnfFFZ5XYIqw94+rnN+Quf0REDhy/5vaHho3+6rbwq8vdzW2nSrSAOMBZZ1vumDwsI6+
EUL7CeNrrFt3MZKWfR08Snxq2F6Q/L4cT8fEYYB6ED84HH9tklx5FY+TGEIR4XZfmV36fS99rhMC
CvzVkoh4x5lJblWXDADWHBWIqZ30JnneBI1loxG/STo5AVC+YzWhxsMN4PwS6YYKL3uzxw0aBzAC
mnG2Kk08cfggm6E5eCD1sy052jmGImFH1ic3DG5WnruFmJs+A9l8G3vJ0vzQXQSJraJVvgiHbv4/
ZXKkJZf0GkSV4yNuruZfvJNnEWy0QtntRUDIMnoIeuOC7iFsUor2haqlhfkB4lt6pX3IkKLZ5pcb
UHr+JCCTW/UBNLYHLRt4E3vO57gwIjb4MWNraowkvZFlNWdeDLdp8LoHVX5V1FEEiyc+AWmrc0+X
a3uWiiv/IGAa5i6W0QtBe2DYanCCZ49Mzrbln31GZAJu4oCyGANtN/V3NYGieWehxLgjGbAcDDKQ
qy+Xz1B4cOmfsc1tdws4lOTyK4AOdZ2s2OCYaXaNJAUx28Rs0RfGL8545t8ULMkbXpp6NgqkCbyB
mtUDK4+kGYyQuoQS3a6D/nKuPde3/Zan4AqZcGe2cdOuN6z3ZytqJXs9cCokdGB2+xsItfGRuKhG
jHMEDHmUyBFskZOdW84c/TS9X4j769S8+rQkRdkJ0rhsA9v6nyJPnasBBURzxpj7hbb13opGsf8s
yPcFqlQXjzMU/IBl/W2RUJkVLZCEz5GiGxZrwD9jIJ95x9QufJz4QflrW0t9zeoPidqj5XZBEIZA
tfQY0B6ujX1cCrIdbhCFN0LQ2nJffV4eR57fJjycXDvv+t9jT5m1tp2xeKghsfaTNP2YhYhS3fIt
xWwxHI7OuzS50XDTaM3dh6ZtPgV/hJbXtlhr72x9R5/qQI6DY2DarRIagkStf4uYCCLS0kC/yd2y
Qiy6hQrE7otd5AwiXjxIRv50BMQCtDqdSMApxCFwJjgp6lNIxT8ev65tmi+gSMGq/9cw4ru2tQJv
AfZK1U+fgONwXqxnmWtbsIZcu9Iyp0My6SS7jibN7YvOT1frm98qTuCXJABubAkFc6+bv43lheRw
jmkm53DbttL5dJ0gueEgR0u8eosJba/8iE3pGA1ysQLzMOmQVSZd+bTYKdKqDM4NHMkjhZSkbdhQ
tmnoIRZT8svlaktcuu4sQB799QxSjQksXzOW7PiXiAIPMGYsVHy2Saql3F3OURZ8YqzQLLTvnycf
ibqRxT09wQGRZ1RTKSO4cnvECZ8tuC3P62BpNPiiT34LFh46TVUeFo/saWaruX+spKuG/mlW77Fu
D0DKBOShrqgM1dp9RRpLXMPSsoLEarQQoCPx2RxJ711jxXw/SkubQMAwrwRo0dm6vs8szJMde8za
VWMtrqbA1fRkVrF7M7zWnDK0uN89WwVfhBfDoN2gJRljdT0kIZ0ipe5iK/jq/C1sP4p0MOL7kZA4
VO99yyM/atSxrD2KxgfxcsW99geh2v6POew/Zt+9pgk2VklGtjVh0WppibJUjULOpga/BggJ6Qps
6cpCUfMQr878hNP1NfgD2CdZ/ayVXXrYDzwfNXGKe/Pp85PuLa29ac2HCwBtcHQt6FiEcL5X/QKe
L94FUVbTUjq4d4S+gTM+Za/7sM3lPrkIxPNg4Jl/FB7RatEsDT8JSbr2vKcGm6rKVHBmaYIBxaSm
Zc7nfSL45GXppRIV3D62MXNTL+uWZcJaV+/f7HJnQ8PtA0qNusc5PyaQGoq6m7Sp7bme31ee04Ef
1879WMUbl8JsQCGaoRi3F13KYsIKB0WjHOXX1Syd7cJOJ64eUTLCCJ3EDJu/GO9JBobqTLNrLNe/
e6wg4AUVMqOaX+U3aXh7e+7MBgxTwTx52cTPdRYcHwNNnklSpxrN9fMUJDKE+HBGoWml5rU7P8Jx
OSGsUUFmJRCD9tM6QgejEahjTbsJK2Rs9YJNhPBD9SJrNeIQym42sdLeLf2rxhLFkmYA1iRRIyi/
qr6tQkl7Jzr0uKOn5jw9tzYDGSy2dJJl6Mqd+qDPum5YMIUJYfbG01yizR6zCBlKkyeKqKE82iFh
aFSaocnU5k6UAl9Y2Gvoh91laHI9IINqa+EdqxMw++RGKzeViODv1HbjeDRoBCgvh2HEv51dMnSb
Qy7CqANHxdFDUDAf5HwyqqUCYPbgoo1BFYN2FkUoST7aMiVs5ZudxuDj+gcOpEYSr4ODfdQrpHY6
7WioSXFHr86nxGD0KDIJ9knL+Jq2Ll0mhXTAZPRwoddJjY58GA3THvHJ02K0Vi8XTU+1j3E+AlcS
HNgf4okwd3Ii6fNk1W1GeoWmvnT+iwZ2gqOoAUXoyYaFDWeyjExpW3NpV9F7MpWAW2BLBRJoMpxb
j6jS3mX2D+dSKBXFNST5wY3qtRkbOKRPLT9/SPgw8Ld1lNWLRy0+ysyRxeguEUL9aCfN/N8bYbhw
Z9TUrFn+kuvTZ7H6zJ5VCdMIA9Ash90RXFg0zIjkJuAlfC6BC6OFnv4DHew8BeL84EwnZbZtUMb8
33cmdIMjD1Bzkv2bS7e18vR8XG+qNy7kjecn4Bj223vx5frCszi1+UCIebD/n/WEuyKZvXyd4Fp3
rm7FGVJAddLYOHC2ZXh12qy9QUgoCUFa5NbW1+R1Rp3BlUWpd8g87d/80V+F2ihUNcXh8qfjkq+s
cFNm1qjBmWYXEb8b/OeAaMd0JUmz1MFF4TihtOJEKo3XatBIiIsb9KaznOunEiyI6x+wRR7HVbFr
4BplkAfR0S3o3EsGqc56MyLn92vJDuSdxfQadCc6Lsl7HRTVt5LUwDkkgFF3bVbOSXxOZFcRvoAA
gBjjeYj16A0BD7IixMSISzYI+ojAfDUylLRAr49ER0tTXK9lDW1s09L/STYClUZZg/4ZXdpCDZC+
bgWpy+w6fvBLG2U+Z0nlTW1DHmhIItfvjOewBNBeRsqJ5aowJy+yUqI+VutR6iDWAQeePyNBVsSc
LQVQ865mbFjh6dZtOGro1zaqk188UVYPE16fPAXXkTJnz3yadxo7Kd8dnAapPOEGK5sheDbfWGTU
VvKbl5iR9qUAk3xc9UckSiR2pBIbfS9G24zOSGsUAOcMj63VuvKzRmWTjuJu1kDpkSQeAiekhsDo
vFYNUX+JMvFLcRlVnZoqokxiBDI0xnK1Icx110hgJliRV3GpMdq+c64EuK0AMOra82HWFGrUbfwi
8yOoqtPAurKK09hAcoMmZl7PB7AbOp3rBbIdL5YydVRF8vrFIPelcmv6OzQTEE0X2RGo4aeJq0XV
/l+CcN+LUPosPllY0+vBPHErhiUhSvVuAHCrrAyTq3PiRuRw1dWZNbG4APIVK4CuaYB7BK5f3UmY
G0l7CiiCU6Ay7zaCvHvucznMO0jEYKwYAkjqottWVWlEgz8ZrfxaCY7nfVNcDEOGAfD9VW+CMSsA
IBBFs4FTkME9fEkqyYfauR5PhNr5Y2ryZ+ugl/TBXVkdjCg36qugqH+ZA2bGnlEgHnIbSqlLv+6H
hig35IdUQzWLCKldJ5cRmUUZxcygNbzfBdpiVu5OctjPGo9LlbrT/3lhsTh3wIosFKip8tQHcP1t
etIgzsR+n194cO2z+VkpRBveiXEc/s5sMgUobUNwoFlV/3E3MbCKOYvvutywKQ1pKlwDzgbYhvV2
iH26DuipcSYB+OWQTx2UkI5237kEW9xBEWS9cTlaMlSBc69TE6YoHL7BLyvqdguS1bXrZrR4Q7G8
VKZ4grgVEnI1e8KybBc5GjF1VFernsc1o+WdKtN3c9GfNRNKnW3983XnGhgzTa56uHO9xiX6XVEc
eFaYrPVCsDMxEaWJtYSZEvh93n280FdEIVDkPgoUzXSg9hJutmt0grl4H3vKk8Ccy6SKkN8odHCV
XRTv26sOwr51f5gcqakJorLCCIxRE+egIlQHE0nFtY32wkNYy3k8eiPBSh/KBlZZtFS8zD8H1U/N
yktzgohN/4p+nFsQabi+Q8DxjeaMP4Bplt0vap74QcXyp2DR10Ux315YU3rUyAJLTT74jwMpZqP/
449htZ+pRwuNbSbs1ks6js23OJd49BMrrF5t/24RBWPlX9dNW6Q6899oNc84PiKbkZF45V62oKd2
4NSbr/eFJYs1+518q/6P9bwrgd00L3ekKeBZN8zdUyXSPWac77V3AAGmhS1mZyDIrODjK1XZ+mRW
pmDdbzOcXjf5NwTtEZBYTgYJj4bSVnXhaPCjLN8o7olZBICwFqOIjq9rA88DiQt5V9reabChaQbX
+XlGG+n43m0Co1DsEEXMP7OsI8wPKY/8I0muO8jEm5k0x4iYLe3CRvzW/I88jNvklAtl4Ym3G7GF
mkr9fsM+e8SDUGSpNRbBqICYPx1SBQk4+xBs/wc07Ndi6utlzPPP3FJginEpJkkufhm207VbtGyV
wG6ytecre/0emFcquFCH9RyoxX3b3UC8hKIv+sQfrybgvKQhvpgVeo5Jw/VBFZB8KiGEnEfSEcN5
F+Hm5me5FLDV/QEXOXycE5iMjYKVHC6hiS3JPckbi9jEWucNxJlixn01UafW612USBWxxsrP8e6W
W+o5VDH6yhUuCwuqszZ2M9Ig8iUZRJbTW0aHfKA4l95bn2U4A3Mo44+lmbURzk5imwRJ8VH3Roja
oK6GSsyNzWeu1A3Lkt/22vRAGSs10UpAlCqEyzC3GUcKYKa6C0BvPypngTz52wW+Yf1LqQXGCLWX
6oYM4CZDZvUewS1RVjswOMR6Y/05eLlGCawkI8dUSLqyEvR2PfIlZ7Bk5ubY0yuQYXxKk1Zb7YQM
2kflTBde7QdS6AhyrEmciRFtv+gxZlGl2TmdTbM521Ft6a/n6cNfrKbP6TkOS0JFBdv4IIQubfUf
lFCNVxOFUZ6cbbcgcwpRfPADnA+59Q7fPCyfciVoUxn4Os2xFVoU3BiQMIVA5RtVlh1SLSuofLhJ
NYLLaopjpmu6H+DKajLq0iAtaF0Mypx1uDAYXhtqPJDKAh665wwVuXeCa2rGl8eT4yvDIiJh9SwT
7y482HB6vJu3gC2CGNA9Dsoijs5bzsz7ai0La3XYHm3AT+hCmkuSLbnwUtbw+dQeqOSPSd/ckk/M
0HZPOgllL0ZbehA6h4/wGppdTEy8BTXsnsQSdDgG3FZbBdO8p7fdtKWkebNJHL9QydbaQML/E0H1
PCU28Lif6DM/kVcYM9G97dNzYGd3dXkZSkMkmPtZGkd9gqtDHV7spW5OaRzgv/oiLK4W9THph5Nl
dOd1GNA6mZ8dLE0GkNSh4h/3pvs50XNto3OulVU2pOLICmrQfGXriCytuJl5M4gvGkq7cRVSjq3i
Ac9z+TDX4zs+3uVg/tUhLWl482ZNsbDyicyMVvBVceCjl7/rRPVk2e51iAnh5woRoXkFOu00cuOt
rqD+Cem/ZYVzfpLyJiGRUyRGVUb4bP6xVO4fCYntuGEM3QwTw2dj83ZFsyRzgMpIzMfulIQpTPTr
Sar05oCc7J95yRvAodhhfS+Cbb46edEvovMdvmaPPcpEb4B491rKLNR9zjwTM1gZlsSuDMMRnqtx
RnS7doJTORQTNS7L1hdifvP1D2GQdD1UMFHLd8iIBmfg+UR4I8HaFsZG6K9hu6i68KcVS4cJcsr1
GSDYXP2fh6nwf/TUin4CM3oybZBQ5P4KJjRltFIH/C/OuWvqvCeRXDZ8g4AicJwMSCjPskAgajuL
JzoJMu+XbFH8vctYQyjTfMKgPwjWaJ/05Pywa7WHvgSrxoMOGLumpDaszrTfTXuBenT61IrJR91p
GKY8b5RvbNi0VG1JvctN/V/PJ5+sSVoQwYhqMIw6VznUT1SSIOT4vBvgNl2EXr29p5jZmmNIjOmo
p050xPFEAG4rs+N5n7WUMnDwCsQg56pQVHRNjXj+1fFZlqSCyNT0sIl6Ns5vPkAJrUe7jneKiw8U
EyVqZmoJU7lKgZbKLR+GaO5aYy9Z4KCjHXt7O3sFAczuu1pkwuIKeJANRdo/HzeHPTkdGmvIB+lG
tcTvXfZslsUEbam2SrVDz0GqZBIwlT45rzOaQsg5+YyWhvHJ8lumhpCkqwXJrBd8Vbe1nbHVDNPH
qmHsrqpwUHQxBDrNNxkBCLHTHgvOl59Zc2pDfSRRUsfWMh4QOeOQnaGpFDLvzmXr8JTWCI1QLDVv
ZKLq09kGawo6oLRBJWWgjdPESbGezvPF8i6xMOylk0c9XtVYWzSXdRK1L0XrY9kBukbCE41tOw6+
FT4njjtqoGXp2BSQaIf5LFsh6J9ZMqh2VSXdrQvpX2kbHmrulPXsRAAtaflzIsZ29JRJ6cxcIjRl
vH30jf40nLh/ZEjJaQhjdhnKwNHLJLQH1lhLHR3IuovmzSQeRSoVkh++P53Vcw20i7fKcDvPkI3O
XHECq0AAbOpV3c1oSzKhi183XYDcZc3yWYuIkVvtMsCnze/5JO/dfcL4zg5XvV64TipgxvY4qorF
HDHun4Hqn1EHPviPYwVHuse3lBhcv+UkqWOb9TsYQYUZZooVruDZPuS6U7YEmdEpz8uI1ySbrU4F
xq7fZe5DGd87NWdXvZfW0a5PeC2WG184yGRVLhRiPAs7vjJB5O/0+hOjc1D5f5rE8CpRbAm393Vz
1YU1C0oJmCvJEtWAfznOiXpBtBezEwH/WU9mrIj07rvA9sHXVnO+Jjrx7hOP+hsNzeqAUSjDTZ/k
nWD80dVOLZoldpUo17zfdfXvb02ebpghuElopNxDL0UhitPA1FjcUDD9gHKcv9ITvFVHswKJmkex
rpKfpj+UWofeHihWj/VhGKCDBp8QCYpOY6CuGpK3j8lHms3CFZtdS0KDAqY5EAjhrhHBUUtJBHUa
C8ACb0w4Rq/gYfi/MEtRMhzBnc1NBonBCggzeJwifpY8yu4xDbF/HdYkP0fD6TujQ6K4I8yqNzop
gBcLrrnZeX5FG/fb1sEOOGzBpAos6K0MwwUmTSUEh/RS3w6u5JVGPd+oTh82Gtcu5D5+afAO09A6
+wq1CUtcd7mwpG7vGSxU32XBSQqRL01yBxIiNc5lUIJgmKvGwrk8X6U8ZXoWj2Zsc6Y4PimKMhUh
sQ4OL3+pQ2mYfQJwtNnP7oqe+Pm8dQ4qEFcC6maXw215Z2Ods35SbPcld2hWj7XXNpY3QzymfAPx
jvBWisxSIO2EDoZXLSKUsPYeraJvSJ46kCQ4XlLuVbW3plFSTxE9MpmBREotSMkDejTvRk3fjauk
PgFno/ryy2ykaAZXNLOhMUSC0zAijla3vOG+5/Y1xiHts7xn8xPtHDTCk/dxLysu1coZBDb7sbLZ
tS0vo30xEe2x/XOZM1zE0wJRyZeV53/HLINhgfF4VsyBGE4onr2awZHn4LP2hXjF8Isk5H6Jtrc3
cJP9BAYbLCPQg3i6lTUlg6CBJopTf/JLNGN6wLccCK17wGIdRGujNW+3M0HD/mYjcBIrFyPm8+sN
xM9E9D9+B2PPDuf6AHufFlDbnBZx1iqOl2oLO9l9HWpbpYczVtbhPe06TnG+twuu42Du67FI1dTc
g0k4ZQI2HK0frKSWFZ2AiAGRS5/j6e2DgLgd/nfZRDkq41U2y9JEe1nAuVVEBOyeUq8+KFf3+6us
xpumBLmuXZPeCXKVBYRkcdSTNloCPG47kDg6tPN8ZsPG8r+kD7Xrpa2DfpcGcY9kegIMwHHcg2zm
xuPGmKc5fYSx+Y0dX4+yIdaBsc7JaXgsABhU7pswGFSgdFff3SKCbk/kK218wKy5C47OwMr5sCRL
fodBRYO39lvlt5CVE8v1b3s+BH+qY3UBDD7gznlPLMm1oESx9O0L8vydky+mpa1wOKtpqn1kbvrM
t35wPIBZvvQt8d+BXvbWyflzU4FonhfMvD+HJPvozzIlSdEPq05YCyp1s0LBghRxutZYSdRstQJY
WmPEItZce4n+138dwJmGT1/3X99I5IVE8o9VX9UEfse2dDoigP1ZQdXpbjc/icQRf27qITt5ZjaI
EDptcgw+NFIXfqhAm6xc0vI3fgcQxbfthwuXeJyOIYV0e7FOXRSw9o5EaTxL7ETfhosxDAWE9vxn
apPAKGTIw3yfy5PM/TTQ4m9BBXA1WaELFzHWYKECoTnx6mehSch0psnROpG3j7eOEIgYUxC5L0Ag
NrMqWDxCnBotA21SJUnnUqsrsUUviu/4gQfoc9w3O1lZELaF+IrV9BmEbW1ngv7cDH6fmmkyMlp4
tjLKzVy4A/g1Ia+ag7ivwSpBSB/obELP5bmZSlUnXQplrQUInHw+vDk3H3I1FcuIGquHzCZWws27
j5Xp4vNP3oV10YCPjSWq2q2fJt5DByfSmYCApIGEL+dbFKP+VHVsogtVF4ua34NQjMIZDNjUFqvn
xA3oaaI/od+3kRWh73mkXN8wGRWQOTHwqPMGYq46cphm4oe3glPSKU1xbcVvZT+4PmxEHjBFfZaL
6kbDSzILarMGoTQiF4F/AMrINvYlbCl6jZxIsCW7ErSNLl6I6c8kiNGsfopHYxW6Y1Vc+5hUNMan
9HJ1VQc/1dfzWGDbVk0y8KM1etZX+wmWWnXa3iQEqsI8iR8YZirjJwFSIEtqu6MuyqMinE8AynDT
rDXTNYYke8CWMKMtEBpdzhFx1L1wRbADSwBzAmpggSqXBB3K6ESpnFGFf19llBF94Kvsh9EWYUsv
pNAer9pCngdi+U37Lt2YQhnnjcVOObXOYAexC2WF712qdm9TiveZ7V/GQfjwuVjJ1Li1aSQ3aUaR
Sr0w6jwToZeO+0HkNtvA5Ar7c8SXD5JqaLHSHcFPIsiYCI7Y1X+kp/FWTFtBXbAh6fKraK3pXJA3
/ZLeTW7UU48l4HHlo/1ViEajLtx7tSldtSAK83NazLhv/n0AojkWSVdQrX8uq2TlojXQf5+HFOBH
IouGXy1e4fgKLCh75qRRXAIpllMf/iwGvIYaH4agFUYGlb9zHchv1Z1SuX1NFQSdICSTBmlUx+a0
87I8Xm1wfyvM7XT68KoYzIaR7sKsB3Fh3hIzMBtzJx5OwWrfvV3huYqoyXEAwpPGCCANg03aQEh1
9jwAGxGpYimv5SmrGYXvOrjTghe9bpp+nxXa8Z3HNQieMmc41MG/FT5BncKwRwq9GFsaLKRcPlC6
UfwByXOUyHndaBNjNLGDs9ZrJhOxP/P6DGXx+VQz1KoAdgv5cd3cIHnXpjA/J+ybHqll/stKe+op
Y0c7vy1GbZu+5K+XjNGnAFVZQc0yd80Hd8+AtkbPtTRGnrmc0mdBmMnGxKXVqIh8YnIiJTlRv6CX
UPih+eYxGvT8VOSvO37l6hkLGHDn+nFmqQPyNKgsJjb8cRq9yu2TGFdgAg4vc2D3GUb6tA+4ACIn
LQ85opxddcroRDTsylv3GMU4gKOFhhy22xjjzdsA4oG2s107EUM1mMzTSdKyp0ZgjLCTyL7vr4f/
q1Bbwxi+crWVe1QJB2ZUpXe8Yn7QYYoLzWzD9MDvmcjVDvOSmhBpgvfDf/oMVdyrwAUl64Zesm1w
XsNArxNMwMaLaCjD82y4r7ASB1X+l897QTDe8Kxub1yukbQ/8iYaRWWeyioYlBtX5aOnBSgTjo5q
4W38P2hNXcSz5LYPKbyX94KSBRvCVLZDl9ymVeDEr5eN/Jsii4OYnJG5su7YUSmWHCtBcuHeIY+l
N94q+Q5g9HuIStMQAcgmawXiBiXC0VtrBp9InRBNRoyz6fZztb8RgMjSuHgdtbxlYg2nsfawD2gL
8sbcJ9vkpNOS2FiKf9n29ZnN6mPBJt6zt1YAQNQ2szjf7b6Ribi7ZAmGQePN/hLM1+z7WbXOBbP0
NkFAZ1T5Nb2xxN+/pvLgmj+JB6qVLO3mGjyf8YbTFf/hbF48WtHtYCnvSpK5CSKcFkygLfmSLvE0
otcBJzMoVII7r6SMlOST0SXk2f3F81SJ+ejCnl5HRjhk88kDgOfHrvmggkDOEvXUW3vrqgo4bV/T
g0bOaVmC/CmU5GFhsr84laQBqJCbQn4ZrccpCJOrTxXnyjJde6NWVJ1fOBTsQmeQJ2dLMqUWjKrB
d0ZaaPsVAe22dXaRjcvImMVpLy2HL7Th7yTg5Wf/kO0lY2LXEffYj/VHeucUmYmPlqUBrPFcok8H
gh9jQK6VBXVgH68mdRORDmKiEq+VzlHe4l819gm6DNXcOhzwMIeZYeh5GzYk5Y/2+6dJsjqZzrBe
K2HkBnkH4dpda5aVsBOuAEVPtNmbp4zbTmsInvhcPG7y1lUcvOsSov19KYJyzIhxL05doW1DcZgr
DGcRFbwe7cDsLvfkyuSMU2A0Kfyll8YLhhgjnZorsU64PcxpOKibNupbW6M01Jyk3SYJel7JpZLp
RcrnKdrCU4X6gAEldjVu4PL2UxJmkvt0I335H9cOtzhL3/nmP6BSysFQParQHzPR8eiZFXaoTg24
CX4+pqG4MNOAnBggRzN2d5NF6nWt3fGzNXGkOYF4vV+t94vIsvWZs6kWApSFmi6kC51trPbJeG7i
OMHuehB+FwLksF2+Cr37CG72X2TE+wkh9hr0YSM680kQ4JOVFDzh0eW8y5xgupfA1NF9P/KJN3A7
qHLudjYbm1ruiXvCHy0HWChcEvZeFKeRzF/vOMJRXOGLv07iisYGQozBzA68LFZETKdKddxmi8sR
62hsZytAeciajCm3vIkkZFJQ+hmit4W8FBpT4RycmXGj4XmTYl4l11D0vjdRx5aAiUeWcPr80z+X
8mw3v5tNGVixzBAo1kWjDmH0XzheDltuOiTClmMq2g0Z47dqib4rawUA+Z8XLlYjSooReIwM9Wah
zFlIfCeHHawAw0/ehjHj7s0LWsN9UrtWKcLYbjhFvd2srYBVIDxhG94if9t+rPQN9MRWzry8QH1q
nzh79zxshIt15DFj204O7xfTDm3YwnUPI2RfShGwF+vj8VB7hmsLoeA41oN6LcewryPGA50WGfLh
5P7GhwGX4zzqrcMTjAEQZXgxLH+S2QPrLCD87xI7s3ijQkoEcaBDyz3L9PTkI6WhwWAY4b4G0Dlr
f3yOmtnWx90o+1ZYJu5Ktr8drk1hoMQDdsrkaX/eTQn9RlRaZi5bfBDbXT189bxRwLLz6u+NBirp
JosMNYSVCz1fhWMJvA4QlrQ+d73A2GgkYXg/GYWdptzCCPabGcR3CIigTfDBGZ3jtOTycNejmR7f
0RJS1QV48LYRa9rjWAM15WCh/nCpSH2SY1eRL7IIpk3qesMC48suwdpWcTM/Ne1e2R1WzlPSh1cW
GhRragiyC5iqEJUWRvKYzUrrudtSJ7NbeaJu7iix5AIohcn4F7vTCVAKjPfxsBmvnIokdpHbxU6w
PtWO343oZ3/2Dtu6fJ9oLu2ILMFwnBtOsZF8GoDf2yf3s3OH8Xl73tpyssGqEiXLoqvTfHKt30lc
m52iEcZVcwanzDab7D+wtbYxKj0cftYNouhrQPLkY+VG2ZBdybqPCmn+bGpTNsWlCECzo9kf/Vu/
vCfDuCnrGIJGgfGnCxXIEgkiylTOuWmnoPu2rua2//bNxp8KF+eGbwOTLhlvZGfx9elDldSmT/Q+
dnN5nrvzp5qeRQvLzPAzmHs+zb1AXcFSPSsXozGsGDQwd3oHnHFXVZsv4iPRYXx7Gw8FBDuQty0c
1Y4M678L3hKbvvjQ7RMv1hEnda0iMk1eJjqbxcppvzroKHfr3FLVcT9ItAyEUVYxxZaMAhALJvYe
uB5JeJB/UIEDE86NNouIH7xzaGqsL3v7c+bP9dZ+ZiYiSeSZrNFDmHXKvUr6W81xz7OmCk0QD/54
2faxMnQF/pzbWQy6hN6SgIdldtlXYnAQhOKK+TryrNcpyCyu25xVc4EywfY/b5dvZyMPQwKdsZy6
eh0jq7cfFrnbcAXclm6SSChRYZVf1DfOxagfvKBS4mpPFV8sk0zdsB2+Bmri3++OilP/M6X9siE9
UAGNumqtShCpOaBpzPcaAllosFT3dazew7bYmyTWiJRjN0t+Ou4GkfznqeG/zaDxMmUkBH0c2i4y
UGDZlB4RG17PJGpOOWcFjsmfWM5XXiupCXZLssnr7oxJCE/XqYxHVBBn18lKqayaYSNbob6fhKmE
oAZb+VwT68qk3bwIjfvxpvoopwgI3bcjmudnWbpPOq5udxO9j2CcGSagheV/+SCPUnzt5N6NxXJ0
MU3gJqlTyRvQ4zwx4gtoHbizNTolwaS1Kw+3x2er/QvLyXZIwdeW+3ZcbqaWO2+Nu6Um4S5H+CzP
w/EySXW4TGFVF56D1uKZxdykQiRpUVELyQkQrtC9sHXGebBt1+BY+swL6FT5CKPDW8BpXCgU7dh1
QGFlaTKRYsFMF5kg9RLZJ7dJRoUwN/5rNm02S767Ma6wj5Ay13joM3fIUzHaUanzZFtxN5dn4tq5
S7Cr2cBuNNzmWLiGAKy1nFt3W7OgB2zjwmNkbD2t2KcBSMUV65uwidUT6lGKNFyA3A6B6olZWOVZ
v0/+LEUTdpc+ifyvAPnuqB/IxG7s8PC27YhbNMVVRvlR3iZSV6PmSILZe6edWthM5Hx7LNbTIRRC
KaS/LnCKhvN0L7fe9NmzdRARBh0aQRAo20ht3cmtb0QVD4SMUrDHImsg2FcXb0o6nBlM9Hs9d19I
T+pnEpZk/ZxagIu+jyHTTfbJvvcoIffGhzabPd4cWtbLkNnvkk6ZYoDc9dMlY7iS210WMSqAX4AI
pwk8ZBUSS30d+LA6IxHJe7lpB+L/V0dqSOFTRv2VNH/ra4AKByl/5gvb3g+bSnjrIsr2r3O9OJ/v
ho/i2TVf+yd5uZ8NRCgoX7NPbuuM3jX77xBxhvYDnLTIKzYnhFfrSsdpEmrbvmXzKUJML91StCYS
OILZYnwjR3eKn7qAz8cX3cDUs0Zw7lt3B1clgcexWE4euilR0ZwtKnGwgbtcsgYsUVJ0Fl05kdhX
9j+d7+YP2X33GbB0tUD9pLzGo+PJ/MCX64/eIaxCwukJ1iXOVVuqPeoubBNBuCPfrIlyxuE7uv0D
Bt+1GILxkdw54rXJ87e/4Lpx2cublXK0v9FKEbnncK249VLKioGryO3zIUyvtPjZqsyNpskpVN+3
pCBgNYi/5XuAZ5xSSmtt8TRIGFl0ynLA+4AwDk4xIFp1YlF+SuCcPTIF4zmr2lV01OGcRCehW6s7
mPgXJrtLu2hptoe3A6bObMcQxcFvTTW9y4qU0Gn8JtDldMq2HSIXXAr9ZcSfG/tegquU2tGFesKV
MH0w3eAO7VndDTDJyz0oxskxVvBjUzfWTwVwEFsIRXdZiDCNNPIgFrkjtqBI9X/XwgbEvDrNx3dF
P7tsFnSOk5v2msti0nAUaf9DUij2T+jp9o/CB8cDJMqSqga1qtm6tzYQ3VddkUaVNnIpzmFqSVc8
x2+DpYKSOTKp+AQCkTHIZJVnI/4WW7eEg3zP91e8B6o3IezenLv7LR+VZZquxRWRahfbEizyYZOA
Tt4ERHQ2qLY0fGoVflSPgaypsP3NU1oaqz7QEuYIVJS2ICotuna3AN+Id2EzHZy2lsg8j3k4fY+h
Ht14Bk1We9Tebw2iYMmU6qoz4YNgmkkT0I8XWjro3B2EmsozlVxxciHPl4P5B0YIhVIkQYCJPX2S
pbihLvRFnYxqWyJP1uBQBiwzi/me93H1TguDILz8bJIGjJULNMu7XKe8o3nY4OdE/sO9AZAi2Z7t
lswr/3vjYqFqsG7JDHdDiXxo4BT/N2Mk2nCrQUz5rBpOdT/HZLPbyTcvO39F87ms9zDUG8+JQiYb
qMXlTPDWBk1RThFh2zbTdaPjvjLnMwcJzYvJB1dVh1UzHeM7zrbQJkZFkMj1E8mIukIHiXZ0giyG
jadO/ezJ9TOzLx4t/blGw2/QvcecXcbpIMP8BIybad4+vFmXFUmNZd6qyOGkVtw9fGLGcrv1jZ8Z
e7lNtsAs8Mo2Jpdq0mr1AsxVHxX9JyVuohGjZYtQrKFwEcY17bXUB2beYcis043UpEj7xC1VlSg4
BEUtlu0aAYH4qnrrBpV1hv+7NEf/m6P+62mY4++JW4ANFRjzb91Va3UT6EE2xNzow7USp6W+iSa/
VrLUR/bNFQa3VTSLJAkifUMvp70+BE0rJzCVE5ZQ1MXamjWKtsuJAsBKYq7ykneaZt8QI2h+a/py
ECaAtu6kXwdtIKSjq3BYAZpgp2BVmseAXS910RJGhrxQjLhy3TCU6ccxeusW0UH5RzewHyWhsb4J
B8wpsVeZY7OD6eCNWSvUl3IMLW4edIbdVexvJNVJqRsA4/InhsR/Ss/JrGYozWflCZiB9Zz7PRkt
sXLeXcY1fSEaqV5kWzktdnz607tUja0RBrbo0TTXScPmz2NnQ2CNHAeSmTODgjEDIVB9/f79a4HP
zmqgL+A2dXl49vG9o9CiTswyh9w9GyMbDA2VwM8uADWdxIqI9eACGaQO6GrbtP88GpRPzyw3m6q4
85wpOZxWmrop95M+SFL7X4LbXbv23GSqVBWoiX3KI3kIc4G/9zanWzQylvmUQE0urQJm1qkswkxx
bb/mVr3E3YqY+z3lZPdCSyLeZdzqnPApTbEMIn6gZL3TTx6Ig66CTKSbjsDg2oFGsCUF+FO5SoKO
ttChB2MPA7kBxRRJy0sZztY/4I5GlmmngvjJ2S5nH8TTQ96gCDUxw3u/LoMQpggdRhPN762joxzH
QnI2DhHPsZi4ccys5XcP+M+ura3z5ssC7DdSevhvW8QDGBCHz+V0kNeoDg3isDx6wr3uTwms7Htb
GMHv3b7O/QrHNq+J4rfwfq1VbW7EHJkoHSESNAgAQpQVWXOwUc0ZNdnr99hP0MRidv2iH4h4rD3Z
WIEWJq7q/gPMRf5vMQT2GmPHS8DrYfUdlDrHhUC0lPY/cXnITAtlrK3In3KseOMQxl+S6ePcAA9g
lWUs8yrSrLqPLk01TboMfOgL/FtdTQ+3+EWhxQaLX0yG3LQO4Wlz56T6cdzOrFrvbpNdHCslvvRJ
rw+I+A2X7cp6k4ACefHoOnL0rX3aym3lR/xNyDXcVqXP19gbztfpBGXfbi5qQcmM+ZX0Hocku8qF
I3e6FL3E8zimLy3lpBOqV2mb5TEb+TrVK0c1R4c7pWRAl10VsJcz+pVe0hWmmdcTEr5NDNNqhrOv
O4ndjMT8eD6Zx6ii13PTvPKBokaap67UJuE3lEYoJg2FcTwbsq4uh7s5kLsOCeIcKTPsnTBUI1p7
NKxGF+kZHtshWKM+vUoigzKhQTZovBmC8T0afz1GCr0KKpwtD4b/5Q9XvznWZ5CYOOLAfiDe6g25
gCYZdSlTwm3demoA6lh5Lto2nMdx7B/3ZA7ena0qJD9Mujm/ufcWkgndCmIvlwisRuIiZihgMV7d
H1YIh4qVAr15fp5lTmqje/jBHl1yaLOTQsVgks1nu3FMYW/QWjr3SOs5Bmz8GlxkTMa9Si5zYDQ5
mMSiJfhYJwIU+XvXLF3vFoKZF5/vgpojhvqzgadVg9XYUDi6SuJk8anOzXmHPFgGj+RaWNJHymKD
MYpbSs5agot1oaDOM3+KyjCrWK1vX72S+vatob5DBk20dLsgUgVC0h6aPdr3lYgI5rA2OD/z8299
2c1bIrZeTbbF1VEy9RDrkWArD2VQSasD4sQjcs93UiOtPjlKHny5tmNH4MBpznvx+f7VR+uSyoHb
F6eK9TuyLGy8w/2mzA4v/97w+RHfhrpykiATpIUL47Nma2Tyvij3JwZVf/PwcQDPUU2YoJEmh+d3
KLTlgsPHVUhYSaBeQu/rzP573oT7iUOiX7fLuMNrszIMkLxNao+PqpDZ4p5xPTNdcAbXZe3LTXF4
TWvObrSRBKTynOTy7Ak6LIPeSLP9JzM9Wp67hZ6Hru8+Of2KMSJcPNUnkybcm6/IPkAd1Hs4hLW8
M4HyQrUyRfmExHFWEJ9CqOdBSjutOpoDpipdZt+W91c4CUYjpEhlcaABmvs3rXOIT+ZDqonuv7FC
jvMeEoD5XFE0Uass6ovzCTXoeIwOGXwkAH/TOYLva9AcGhbc59QZzPhgy0qIiAz1E/h1i/xoKnyn
G8OxXS6+mvIWw/nqBMX0H0k=
`protect end_protected
